module mnist_rf_pipeline (
    input wire clk,
    input wire reset,
    input wire [783:0] image,
    output wire [3:0] result
);

reg [783:0] input_data[9:0];
wire [9:0] tree_result_index[9:0];

wire [3:0] count[9:0];
wire [3:0] winner_0vs1;
wire [3:0] winner_2vs3;
wire [3:0] winner_4vs5;
wire [3:0] winner_6vs7;
wire [3:0] winner_8vs9;
wire [3:0] winner_01vs23;
wire [3:0] winner_45vs67;
wire [3:0] winner_0123vs4567;

wire [10:0] next_feature_0[8:0];
wire [10:0] next_feature_1[8:0];
wire [10:0] next_feature_2[8:0];
wire [10:0] next_feature_3[8:0];
wire [10:0] next_feature_4[8:0];
wire [10:0] next_feature_5[8:0];
wire [10:0] next_feature_6[8:0];
wire [10:0] next_feature_7[8:0];
wire [10:0] next_feature_8[8:0];
wire [10:0] next_feature_9[8:0];

wire [9:0] feature_index_0[1022:0];
wire [9:0] feature_index_1[1022:0];
wire [9:0] feature_index_2[1022:0];
wire [9:0] feature_index_3[1022:0];
wire [9:0] feature_index_4[1022:0];
wire [9:0] feature_index_5[1022:0];
wire [9:0] feature_index_6[1022:0];
wire [9:0] feature_index_7[1022:0];
wire [9:0] feature_index_8[1022:0];
wire [9:0] feature_index_9[1022:0];
wire [9:0] label_0[1023:0];
wire [9:0] label_1[1023:0];
wire [9:0] label_2[1023:0];
wire [9:0] label_3[1023:0];
wire [9:0] label_4[1023:0];
wire [9:0] label_5[1023:0];
wire [9:0] label_6[1023:0];
wire [9:0] label_7[1023:0];
wire [9:0] label_8[1023:0];
wire [9:0] label_9[1023:0];


assign count[0] = {3'd0, label_0[tree_result_index[0]][0]} + {3'd0, label_1[tree_result_index[1]][0]} + {3'd0, label_2[tree_result_index[2]][0]}
                + {3'd0, label_3[tree_result_index[3]][0]} + {3'd0, label_4[tree_result_index[4]][0]} + {3'd0, label_5[tree_result_index[5]][0]}
                + {3'd0, label_6[tree_result_index[6]][0]} + {3'd0, label_7[tree_result_index[7]][0]} + {3'd0, label_8[tree_result_index[8]][0]}
                + {3'd0, label_9[tree_result_index[9]][0]};
assign count[1] = {3'd0, label_0[tree_result_index[0]][1]} + {3'd0, label_1[tree_result_index[1]][1]} + {3'd0, label_2[tree_result_index[2]][1]}
                + {3'd0, label_3[tree_result_index[3]][1]} + {3'd0, label_4[tree_result_index[4]][1]} + {3'd0, label_5[tree_result_index[5]][1]}
                + {3'd0, label_6[tree_result_index[6]][1]} + {3'd0, label_7[tree_result_index[7]][1]} + {3'd0, label_8[tree_result_index[8]][1]}
                + {3'd0, label_9[tree_result_index[9]][1]};
assign count[2] = {3'd0, label_0[tree_result_index[0]][2]} + {3'd0, label_1[tree_result_index[1]][2]} + {3'd0, label_2[tree_result_index[2]][2]}
                + {3'd0, label_3[tree_result_index[3]][2]} + {3'd0, label_4[tree_result_index[4]][2]} + {3'd0, label_5[tree_result_index[5]][2]}
                + {3'd0, label_6[tree_result_index[6]][2]} + {3'd0, label_7[tree_result_index[7]][2]} + {3'd0, label_8[tree_result_index[8]][2]}
                + {3'd0, label_9[tree_result_index[9]][2]};
assign count[3] = {3'd0, label_0[tree_result_index[0]][3]} + {3'd0, label_1[tree_result_index[1]][3]} + {3'd0, label_2[tree_result_index[2]][3]}
                + {3'd0, label_3[tree_result_index[3]][3]} + {3'd0, label_4[tree_result_index[4]][3]} + {3'd0, label_5[tree_result_index[5]][3]}
                + {3'd0, label_6[tree_result_index[6]][3]} + {3'd0, label_7[tree_result_index[7]][3]} + {3'd0, label_8[tree_result_index[8]][3]}
                + {3'd0, label_9[tree_result_index[9]][3]};
assign count[4] = {3'd0, label_0[tree_result_index[0]][4]} + {3'd0, label_1[tree_result_index[1]][4]} + {3'd0, label_2[tree_result_index[2]][4]}
                + {3'd0, label_3[tree_result_index[3]][4]} + {3'd0, label_4[tree_result_index[4]][4]} + {3'd0, label_5[tree_result_index[5]][4]}
                + {3'd0, label_6[tree_result_index[6]][4]} + {3'd0, label_7[tree_result_index[7]][4]} + {3'd0, label_8[tree_result_index[8]][4]}
                + {3'd0, label_9[tree_result_index[9]][4]};
assign count[5] = {3'd0, label_0[tree_result_index[0]][5]} + {3'd0, label_1[tree_result_index[1]][5]} + {3'd0, label_2[tree_result_index[2]][5]}
                + {3'd0, label_3[tree_result_index[3]][5]} + {3'd0, label_4[tree_result_index[4]][5]} + {3'd0, label_5[tree_result_index[5]][5]}
                + {3'd0, label_6[tree_result_index[6]][5]} + {3'd0, label_7[tree_result_index[7]][5]} + {3'd0, label_8[tree_result_index[8]][5]}
                + {3'd0, label_9[tree_result_index[9]][5]};
assign count[6] = {3'd0, label_0[tree_result_index[0]][6]} + {3'd0, label_1[tree_result_index[1]][6]} + {3'd0, label_2[tree_result_index[2]][6]}
                + {3'd0, label_3[tree_result_index[3]][6]} + {3'd0, label_4[tree_result_index[4]][6]} + {3'd0, label_5[tree_result_index[5]][6]}
                + {3'd0, label_6[tree_result_index[6]][6]} + {3'd0, label_7[tree_result_index[7]][6]} + {3'd0, label_8[tree_result_index[8]][6]}
                + {3'd0, label_9[tree_result_index[9]][6]};
assign count[7] = {3'd0, label_0[tree_result_index[0]][7]} + {3'd0, label_1[tree_result_index[1]][7]} + {3'd0, label_2[tree_result_index[2]][7]}
                + {3'd0, label_3[tree_result_index[3]][7]} + {3'd0, label_4[tree_result_index[4]][7]} + {3'd0, label_5[tree_result_index[5]][7]}
                + {3'd0, label_6[tree_result_index[6]][7]} + {3'd0, label_7[tree_result_index[7]][7]} + {3'd0, label_8[tree_result_index[8]][7]}
                + {3'd0, label_9[tree_result_index[9]][7]};
assign count[8] = {3'd0, label_0[tree_result_index[0]][8]} + {3'd0, label_1[tree_result_index[1]][8]} + {3'd0, label_2[tree_result_index[2]][8]}
                + {3'd0, label_3[tree_result_index[3]][8]} + {3'd0, label_4[tree_result_index[4]][8]} + {3'd0, label_5[tree_result_index[5]][8]}
                + {3'd0, label_6[tree_result_index[6]][8]} + {3'd0, label_7[tree_result_index[7]][8]} + {3'd0, label_8[tree_result_index[8]][8]}
                + {3'd0, label_9[tree_result_index[9]][8]};
assign count[9] = {3'd0, label_0[tree_result_index[0]][9]} + {3'd0, label_1[tree_result_index[1]][9]} + {3'd0, label_2[tree_result_index[2]][9]}
                + {3'd0, label_3[tree_result_index[3]][9]} + {3'd0, label_4[tree_result_index[4]][9]} + {3'd0, label_5[tree_result_index[5]][9]}
                + {3'd0, label_6[tree_result_index[6]][9]} + {3'd0, label_7[tree_result_index[7]][9]} + {3'd0, label_8[tree_result_index[8]][9]}
                + {3'd0, label_9[tree_result_index[9]][9]};

assign winner_0vs1 = count[0] > count[1] ? 4'd0 : 4'd1;
assign winner_2vs3 = count[2] > count[3] ? 4'd2 : 4'd3;
assign winner_4vs5 = count[4] > count[5] ? 4'd4 : 4'd5;
assign winner_6vs7 = count[6] > count[7] ? 4'd6 : 4'd7;
assign winner_8vs9 = count[8] > count[9] ? 4'd0 : 4'd1;
assign winner_01vs23 = count[winner_2vs3] > count[winner_0vs1] ? winner_2vs3 : winner_0vs1;
assign winner_45vs67 = count[winner_6vs7] > count[winner_4vs5] ? winner_6vs7 : winner_4vs5;
assign winner_0123vs4567 = count[winner_45vs67] > count[winner_01vs23] ? winner_45vs67 : winner_01vs23;
assign result = count[winner_8vs9] > count[winner_0123vs4567] ? winner_8vs9 : winner_0123vs4567;


always @(posedge clk) begin
    input_data[0] <= image;
    input_data[1] <= input_data[0];
    input_data[2] <= input_data[1];
    input_data[3] <= input_data[2];
    input_data[4] <= input_data[3];
    input_data[5] <= input_data[4];
    input_data[6] <= input_data[5];
    input_data[7] <= input_data[6];
    input_data[8] <= input_data[7];
    input_data[9] <= input_data[8];
end

tree tree0(clk, reset,
    input_data[0][feature_index_0[0]],
    input_data[1][feature_index_0[next_feature_0[0]]], input_data[2][feature_index_0[next_feature_0[1]]],
    input_data[3][feature_index_0[next_feature_0[2]]], input_data[4][feature_index_0[next_feature_0[3]]],
    input_data[5][feature_index_0[next_feature_0[4]]], input_data[6][feature_index_0[next_feature_0[5]]],
    input_data[7][feature_index_0[next_feature_0[6]]], input_data[8][feature_index_0[next_feature_0[7]]], input_data[9][feature_index_0[next_feature_0[8]]],
    next_feature_0[0], next_feature_0[1], next_feature_0[2], next_feature_0[3],
    next_feature_0[4], next_feature_0[5], next_feature_0[6], next_feature_0[7], next_feature_0[8],
    tree_result_index[0]
);
tree tree1(clk, reset,
    input_data[0][feature_index_1[0]],
    input_data[1][feature_index_1[next_feature_1[0]]], input_data[2][feature_index_1[next_feature_1[1]]],
    input_data[3][feature_index_1[next_feature_1[2]]], input_data[4][feature_index_1[next_feature_1[3]]],
    input_data[5][feature_index_1[next_feature_1[4]]], input_data[6][feature_index_1[next_feature_1[5]]],
    input_data[7][feature_index_1[next_feature_1[6]]], input_data[8][feature_index_1[next_feature_1[7]]], input_data[9][feature_index_1[next_feature_1[8]]],
    next_feature_1[0], next_feature_1[1], next_feature_1[2], next_feature_1[3],
    next_feature_1[4], next_feature_1[5], next_feature_1[6], next_feature_1[7], next_feature_1[8],
    tree_result_index[1]
);
tree tree2(clk, reset,
    input_data[0][feature_index_2[0]],
    input_data[1][feature_index_2[next_feature_2[0]]], input_data[2][feature_index_2[next_feature_2[1]]],
    input_data[3][feature_index_2[next_feature_2[2]]], input_data[4][feature_index_2[next_feature_2[3]]],
    input_data[5][feature_index_2[next_feature_2[4]]], input_data[6][feature_index_2[next_feature_2[5]]],
    input_data[7][feature_index_2[next_feature_2[6]]], input_data[8][feature_index_2[next_feature_2[7]]], input_data[9][feature_index_2[next_feature_2[8]]],
    next_feature_2[0], next_feature_2[1], next_feature_2[2], next_feature_2[3],
    next_feature_2[4], next_feature_2[5], next_feature_2[6], next_feature_2[7], next_feature_2[8],
    tree_result_index[2]
);
tree tree3(clk, reset,
    input_data[0][feature_index_3[0]],
    input_data[1][feature_index_3[next_feature_3[0]]], input_data[2][feature_index_3[next_feature_3[1]]],
    input_data[3][feature_index_3[next_feature_3[2]]], input_data[4][feature_index_3[next_feature_3[3]]],
    input_data[5][feature_index_3[next_feature_3[4]]], input_data[6][feature_index_3[next_feature_3[5]]],
    input_data[7][feature_index_3[next_feature_3[6]]], input_data[8][feature_index_3[next_feature_3[7]]], input_data[9][feature_index_3[next_feature_3[8]]],
    next_feature_3[0], next_feature_3[1], next_feature_3[2], next_feature_3[3],
    next_feature_3[4], next_feature_3[5], next_feature_3[6], next_feature_3[7], next_feature_3[8],
    tree_result_index[3]
);
tree tree4(clk, reset,
    input_data[0][feature_index_4[0]],
    input_data[1][feature_index_4[next_feature_4[0]]], input_data[2][feature_index_4[next_feature_4[1]]],
    input_data[3][feature_index_4[next_feature_4[2]]], input_data[4][feature_index_4[next_feature_4[3]]],
    input_data[5][feature_index_4[next_feature_4[4]]], input_data[6][feature_index_4[next_feature_4[5]]],
    input_data[7][feature_index_4[next_feature_4[6]]], input_data[8][feature_index_4[next_feature_4[7]]], input_data[9][feature_index_4[next_feature_4[8]]],
    next_feature_4[0], next_feature_4[1], next_feature_4[2], next_feature_4[3],
    next_feature_4[4], next_feature_4[5], next_feature_4[6], next_feature_4[7], next_feature_4[8],
    tree_result_index[4]
);
tree tree5(clk, reset,
    input_data[0][feature_index_5[0]],
    input_data[1][feature_index_5[next_feature_5[0]]], input_data[2][feature_index_5[next_feature_5[1]]],
    input_data[3][feature_index_5[next_feature_5[2]]], input_data[4][feature_index_5[next_feature_5[3]]],
    input_data[5][feature_index_5[next_feature_5[4]]], input_data[6][feature_index_5[next_feature_5[5]]],
    input_data[7][feature_index_5[next_feature_5[6]]], input_data[8][feature_index_5[next_feature_5[7]]], input_data[9][feature_index_5[next_feature_5[8]]],
    next_feature_5[0], next_feature_5[1], next_feature_5[2], next_feature_5[3],
    next_feature_5[4], next_feature_5[5], next_feature_5[6], next_feature_5[7], next_feature_5[8],
    tree_result_index[5]
);
tree tree6(clk, reset,
    input_data[0][feature_index_6[0]],
    input_data[1][feature_index_6[next_feature_6[0]]], input_data[2][feature_index_6[next_feature_6[1]]],
    input_data[3][feature_index_6[next_feature_6[2]]], input_data[4][feature_index_6[next_feature_6[3]]],
    input_data[5][feature_index_6[next_feature_6[4]]], input_data[6][feature_index_6[next_feature_6[5]]],
    input_data[7][feature_index_6[next_feature_6[6]]], input_data[8][feature_index_6[next_feature_6[7]]], input_data[9][feature_index_6[next_feature_6[8]]],
    next_feature_6[0], next_feature_6[1], next_feature_6[2], next_feature_6[3],
    next_feature_6[4], next_feature_6[5], next_feature_6[6], next_feature_6[7], next_feature_6[8],
    tree_result_index[6]
);
tree tree7(clk, reset,
    input_data[0][feature_index_7[0]],
    input_data[1][feature_index_7[next_feature_7[0]]], input_data[2][feature_index_7[next_feature_7[1]]],
    input_data[3][feature_index_7[next_feature_7[2]]], input_data[4][feature_index_7[next_feature_7[3]]],
    input_data[5][feature_index_7[next_feature_7[4]]], input_data[6][feature_index_7[next_feature_7[5]]],
    input_data[7][feature_index_7[next_feature_7[6]]], input_data[8][feature_index_7[next_feature_7[7]]], input_data[9][feature_index_7[next_feature_7[8]]],
    next_feature_7[0], next_feature_7[1], next_feature_7[2], next_feature_7[3],
    next_feature_7[4], next_feature_7[5], next_feature_7[6], next_feature_7[7], next_feature_7[8],
    tree_result_index[7]
);
tree tree8(clk, reset,
    input_data[0][feature_index_8[0]],
    input_data[1][feature_index_8[next_feature_8[0]]], input_data[2][feature_index_8[next_feature_8[1]]],
    input_data[3][feature_index_8[next_feature_8[2]]], input_data[4][feature_index_8[next_feature_8[3]]],
    input_data[5][feature_index_8[next_feature_8[4]]], input_data[6][feature_index_8[next_feature_8[5]]],
    input_data[7][feature_index_8[next_feature_8[6]]], input_data[8][feature_index_8[next_feature_8[7]]], input_data[9][feature_index_8[next_feature_8[8]]],
    next_feature_8[0], next_feature_8[1], next_feature_8[2], next_feature_8[3],
    next_feature_8[4], next_feature_8[5], next_feature_8[6], next_feature_8[7], next_feature_8[8],
    tree_result_index[8]
);
tree tree9(clk, reset,
    input_data[0][feature_index_9[0]],
    input_data[1][feature_index_9[next_feature_9[0]]], input_data[2][feature_index_9[next_feature_9[1]]],
    input_data[3][feature_index_9[next_feature_9[2]]], input_data[4][feature_index_9[next_feature_9[3]]],
    input_data[5][feature_index_9[next_feature_9[4]]], input_data[6][feature_index_9[next_feature_9[5]]],
    input_data[7][feature_index_9[next_feature_9[6]]], input_data[8][feature_index_9[next_feature_9[7]]], input_data[9][feature_index_9[next_feature_9[8]]],
    next_feature_9[0], next_feature_9[1], next_feature_9[2], next_feature_9[3],
    next_feature_9[4], next_feature_9[5], next_feature_9[6], next_feature_9[7], next_feature_9[8],
    tree_result_index[9]
);

assign label_0[0] = 10'b0000000010;
assign label_0[1] = 10'b0000001000;
assign label_0[2] = 10'b0010000000;
assign label_0[3] = 10'b0000000001;
assign label_0[4] = 10'b0010000000;
assign label_0[5] = 10'b0000000001;
assign label_0[6] = 10'b0000000001;
assign label_0[7] = 10'b0000000100;
assign label_0[8] = 10'b0000000100;
assign label_0[9] = 10'b0000001000;
assign label_0[10] = 10'b0010000000;
assign label_0[11] = 10'b0000100000;
assign label_0[12] = 10'b0000001000;
assign label_0[13] = 10'b0000001000;
assign label_0[14] = 10'b0000100000;
assign label_0[15] = 10'b0000001000;
assign label_0[16] = 10'b0000000010;
assign label_0[17] = 10'b0001000000;
assign label_0[18] = 10'b0010000000;
assign label_0[19] = 10'b0100000000;
assign label_0[20] = 10'b0000000100;
assign label_0[21] = 10'b0100000000;
assign label_0[22] = 10'b0100000000;
assign label_0[23] = 10'b0000000010;
assign label_0[24] = 10'b0000000100;
assign label_0[25] = 10'b0000000010;
assign label_0[26] = 10'b0000000100;
assign label_0[27] = 10'b0000000100;
assign label_0[28] = 10'b0000001000;
assign label_0[29] = 10'b0100000000;
assign label_0[30] = 10'b0100000000;
assign label_0[31] = 10'b0000000010;
assign label_0[32] = 10'b0010000000;
assign label_0[33] = 10'b0000010000;
assign label_0[34] = 10'b0010000000;
assign label_0[35] = 10'b0000000100;
assign label_0[36] = 10'b0000000010;
assign label_0[37] = 10'b0000001000;
assign label_0[38] = 10'b0010000000;
assign label_0[39] = 10'b0010000000;
assign label_0[40] = 10'b1000000000;
assign label_0[41] = 10'b0000010000;
assign label_0[42] = 10'b0100000000;
assign label_0[43] = 10'b0000001000;
assign label_0[44] = 10'b0010000000;
assign label_0[45] = 10'b0000010000;
assign label_0[46] = 10'b0000001000;
assign label_0[47] = 10'b0100000000;
assign label_0[48] = 10'b0000001000;
assign label_0[49] = 10'b0000100000;
assign label_0[50] = 10'b0000100000;
assign label_0[51] = 10'b0100000000;
assign label_0[52] = 10'b0100000000;
assign label_0[53] = 10'b0000000010;
assign label_0[54] = 10'b0000000100;
assign label_0[55] = 10'b0100000000;
assign label_0[56] = 10'b0000001000;
assign label_0[57] = 10'b0001000000;
assign label_0[58] = 10'b0000001000;
assign label_0[59] = 10'b0000001000;
assign label_0[60] = 10'b0000000001;
assign label_0[61] = 10'b0000000001;
assign label_0[62] = 10'b0000000001;
assign label_0[63] = 10'b0000001000;
assign label_0[64] = 10'b0000010000;
assign label_0[65] = 10'b0000010000;
assign label_0[66] = 10'b0000000100;
assign label_0[67] = 10'b0000100000;
assign label_0[68] = 10'b0010000000;
assign label_0[69] = 10'b0000010000;
assign label_0[70] = 10'b0000010000;
assign label_0[71] = 10'b0001000000;
assign label_0[72] = 10'b0000010000;
assign label_0[73] = 10'b0000100000;
assign label_0[74] = 10'b1000000000;
assign label_0[75] = 10'b1000000000;
assign label_0[76] = 10'b0010000000;
assign label_0[77] = 10'b1000000000;
assign label_0[78] = 10'b0100000000;
assign label_0[79] = 10'b0100000000;
assign label_0[80] = 10'b0000100000;
assign label_0[81] = 10'b0000100000;
assign label_0[82] = 10'b0000100000;
assign label_0[83] = 10'b0000100000;
assign label_0[84] = 10'b0000000100;
assign label_0[85] = 10'b0100000000;
assign label_0[86] = 10'b0000001000;
assign label_0[87] = 10'b0000100000;
assign label_0[88] = 10'b0000000100;
assign label_0[89] = 10'b0000000100;
assign label_0[90] = 10'b0000000001;
assign label_0[91] = 10'b0000100000;
assign label_0[92] = 10'b0000100000;
assign label_0[93] = 10'b0000000100;
assign label_0[94] = 10'b0000000001;
assign label_0[95] = 10'b0000001000;
assign label_0[96] = 10'b0000000100;
assign label_0[97] = 10'b0000000100;
assign label_0[98] = 10'b0001000000;
assign label_0[99] = 10'b0000010000;
assign label_0[100] = 10'b0000010000;
assign label_0[101] = 10'b0000010000;
assign label_0[102] = 10'b0001000000;
assign label_0[103] = 10'b0001000000;
assign label_0[104] = 10'b0000000100;
assign label_0[105] = 10'b0000000100;
assign label_0[106] = 10'b0000000100;
assign label_0[107] = 10'b0000000100;
assign label_0[108] = 10'b0000000100;
assign label_0[109] = 10'b0000000100;
assign label_0[110] = 10'b0000000100;
assign label_0[111] = 10'b0000000100;
assign label_0[112] = 10'b0000000100;
assign label_0[113] = 10'b0000000100;
assign label_0[114] = 10'b0000000100;
assign label_0[115] = 10'b0000000100;
assign label_0[116] = 10'b0000000100;
assign label_0[117] = 10'b0000000100;
assign label_0[118] = 10'b0000000100;
assign label_0[119] = 10'b0000000100;
assign label_0[120] = 10'b0000001000;
assign label_0[121] = 10'b0000001000;
assign label_0[122] = 10'b0000001000;
assign label_0[123] = 10'b0000001000;
assign label_0[124] = 10'b0000001000;
assign label_0[125] = 10'b0000001000;
assign label_0[126] = 10'b0000001000;
assign label_0[127] = 10'b0000001000;
assign label_0[128] = 10'b0010000000;
assign label_0[129] = 10'b1000000000;
assign label_0[130] = 10'b0010000000;
assign label_0[131] = 10'b0000000100;
assign label_0[132] = 10'b1000000000;
assign label_0[133] = 10'b0000010000;
assign label_0[134] = 10'b0000010000;
assign label_0[135] = 10'b1000000000;
assign label_0[136] = 10'b0000000010;
assign label_0[137] = 10'b0010000000;
assign label_0[138] = 10'b0010000000;
assign label_0[139] = 10'b0000000100;
assign label_0[140] = 10'b0010000000;
assign label_0[141] = 10'b0000001000;
assign label_0[142] = 10'b0000100000;
assign label_0[143] = 10'b1000000000;
assign label_0[144] = 10'b0000000001;
assign label_0[145] = 10'b0000100000;
assign label_0[146] = 10'b0000000001;
assign label_0[147] = 10'b0010000000;
assign label_0[148] = 10'b0000000010;
assign label_0[149] = 10'b0000100000;
assign label_0[150] = 10'b0001000000;
assign label_0[151] = 10'b0000000001;
assign label_0[152] = 10'b0000100000;
assign label_0[153] = 10'b0000100000;
assign label_0[154] = 10'b0000001000;
assign label_0[155] = 10'b0000001000;
assign label_0[156] = 10'b0000001000;
assign label_0[157] = 10'b0000001000;
assign label_0[158] = 10'b0000000001;
assign label_0[159] = 10'b0100000000;
assign label_0[160] = 10'b0010000000;
assign label_0[161] = 10'b0010000000;
assign label_0[162] = 10'b0100000000;
assign label_0[163] = 10'b0000000010;
assign label_0[164] = 10'b0000000100;
assign label_0[165] = 10'b0000000100;
assign label_0[166] = 10'b0010000000;
assign label_0[167] = 10'b0010000000;
assign label_0[168] = 10'b0000010000;
assign label_0[169] = 10'b1000000000;
assign label_0[170] = 10'b0000000100;
assign label_0[171] = 10'b1000000000;
assign label_0[172] = 10'b0000010000;
assign label_0[173] = 10'b0000010000;
assign label_0[174] = 10'b0000100000;
assign label_0[175] = 10'b0000000001;
assign label_0[176] = 10'b0000010000;
assign label_0[177] = 10'b1000000000;
assign label_0[178] = 10'b0010000000;
assign label_0[179] = 10'b1000000000;
assign label_0[180] = 10'b0001000000;
assign label_0[181] = 10'b0001000000;
assign label_0[182] = 10'b0001000000;
assign label_0[183] = 10'b0001000000;
assign label_0[184] = 10'b0000010000;
assign label_0[185] = 10'b0000010000;
assign label_0[186] = 10'b0001000000;
assign label_0[187] = 10'b0000010000;
assign label_0[188] = 10'b0000010000;
assign label_0[189] = 10'b1000000000;
assign label_0[190] = 10'b0000010000;
assign label_0[191] = 10'b1000000000;
assign label_0[192] = 10'b0000100000;
assign label_0[193] = 10'b0000001000;
assign label_0[194] = 10'b0000000001;
assign label_0[195] = 10'b0000100000;
assign label_0[196] = 10'b0000000100;
assign label_0[197] = 10'b0000000010;
assign label_0[198] = 10'b0000000010;
assign label_0[199] = 10'b0100000000;
assign label_0[200] = 10'b0000100000;
assign label_0[201] = 10'b0000100000;
assign label_0[202] = 10'b0000100000;
assign label_0[203] = 10'b0000100000;
assign label_0[204] = 10'b0100000000;
assign label_0[205] = 10'b0000001000;
assign label_0[206] = 10'b0000001000;
assign label_0[207] = 10'b0100000000;
assign label_0[208] = 10'b0000000100;
assign label_0[209] = 10'b0000000100;
assign label_0[210] = 10'b0001000000;
assign label_0[211] = 10'b0000000001;
assign label_0[212] = 10'b0000000001;
assign label_0[213] = 10'b0000000001;
assign label_0[214] = 10'b0000001000;
assign label_0[215] = 10'b0000001000;
assign label_0[216] = 10'b0000100000;
assign label_0[217] = 10'b1000000000;
assign label_0[218] = 10'b0000010000;
assign label_0[219] = 10'b0001000000;
assign label_0[220] = 10'b0001000000;
assign label_0[221] = 10'b0000010000;
assign label_0[222] = 10'b0000000100;
assign label_0[223] = 10'b0100000000;
assign label_0[224] = 10'b0100000000;
assign label_0[225] = 10'b1000000000;
assign label_0[226] = 10'b0000000001;
assign label_0[227] = 10'b0000001000;
assign label_0[228] = 10'b0000001000;
assign label_0[229] = 10'b0000100000;
assign label_0[230] = 10'b0000001000;
assign label_0[231] = 10'b0000001000;
assign label_0[232] = 10'b0000000001;
assign label_0[233] = 10'b0000100000;
assign label_0[234] = 10'b0000000001;
assign label_0[235] = 10'b0000001000;
assign label_0[236] = 10'b0000001000;
assign label_0[237] = 10'b0000000001;
assign label_0[238] = 10'b0000001000;
assign label_0[239] = 10'b0000000100;
assign label_0[240] = 10'b0000001000;
assign label_0[241] = 10'b0000000100;
assign label_0[242] = 10'b0000000100;
assign label_0[243] = 10'b0000000100;
assign label_0[244] = 10'b0000010000;
assign label_0[245] = 10'b1000000000;
assign label_0[246] = 10'b0000000100;
assign label_0[247] = 10'b0000000001;
assign label_0[248] = 10'b0000000100;
assign label_0[249] = 10'b0000000100;
assign label_0[250] = 10'b0100000000;
assign label_0[251] = 10'b0100000000;
assign label_0[252] = 10'b0000000100;
assign label_0[253] = 10'b0000000100;
assign label_0[254] = 10'b0000000100;
assign label_0[255] = 10'b0000000100;
assign label_0[256] = 10'b0000100000;
assign label_0[257] = 10'b0000010000;
assign label_0[258] = 10'b0000010000;
assign label_0[259] = 10'b0000010000;
assign label_0[260] = 10'b0001000000;
assign label_0[261] = 10'b0000010000;
assign label_0[262] = 10'b0000010000;
assign label_0[263] = 10'b0000001000;
assign label_0[264] = 10'b0001000000;
assign label_0[265] = 10'b0000000100;
assign label_0[266] = 10'b0000000100;
assign label_0[267] = 10'b0000000100;
assign label_0[268] = 10'b0000000100;
assign label_0[269] = 10'b0000000100;
assign label_0[270] = 10'b0000001000;
assign label_0[271] = 10'b0000000100;
assign label_0[272] = 10'b0000010000;
assign label_0[273] = 10'b1000000000;
assign label_0[274] = 10'b0000010000;
assign label_0[275] = 10'b1000000000;
assign label_0[276] = 10'b0000001000;
assign label_0[277] = 10'b0000100000;
assign label_0[278] = 10'b0000100000;
assign label_0[279] = 10'b0000001000;
assign label_0[280] = 10'b0100000000;
assign label_0[281] = 10'b0100000000;
assign label_0[282] = 10'b0000100000;
assign label_0[283] = 10'b0001000000;
assign label_0[284] = 10'b0001000000;
assign label_0[285] = 10'b0001000000;
assign label_0[286] = 10'b0000000100;
assign label_0[287] = 10'b0000000100;
assign label_0[288] = 10'b0001000000;
assign label_0[289] = 10'b0001000000;
assign label_0[290] = 10'b0001000000;
assign label_0[291] = 10'b0001000000;
assign label_0[292] = 10'b0001000000;
assign label_0[293] = 10'b0001000000;
assign label_0[294] = 10'b0001000000;
assign label_0[295] = 10'b0001000000;
assign label_0[296] = 10'b0001000000;
assign label_0[297] = 10'b0001000000;
assign label_0[298] = 10'b0001000000;
assign label_0[299] = 10'b0001000000;
assign label_0[300] = 10'b0001000000;
assign label_0[301] = 10'b0001000000;
assign label_0[302] = 10'b0001000000;
assign label_0[303] = 10'b0001000000;
assign label_0[304] = 10'b0001000000;
assign label_0[305] = 10'b0001000000;
assign label_0[306] = 10'b0001000000;
assign label_0[307] = 10'b0001000000;
assign label_0[308] = 10'b0001000000;
assign label_0[309] = 10'b0001000000;
assign label_0[310] = 10'b0001000000;
assign label_0[311] = 10'b0001000000;
assign label_0[312] = 10'b0001000000;
assign label_0[313] = 10'b0001000000;
assign label_0[314] = 10'b0001000000;
assign label_0[315] = 10'b0001000000;
assign label_0[316] = 10'b0001000000;
assign label_0[317] = 10'b0001000000;
assign label_0[318] = 10'b0001000000;
assign label_0[319] = 10'b0001000000;
assign label_0[320] = 10'b0000010000;
assign label_0[321] = 10'b0001000000;
assign label_0[322] = 10'b0000000010;
assign label_0[323] = 10'b1000000000;
assign label_0[324] = 10'b0000100000;
assign label_0[325] = 10'b0000100000;
assign label_0[326] = 10'b0000100000;
assign label_0[327] = 10'b0000001000;
assign label_0[328] = 10'b0001000000;
assign label_0[329] = 10'b0001000000;
assign label_0[330] = 10'b0001000000;
assign label_0[331] = 10'b0000000100;
assign label_0[332] = 10'b0100000000;
assign label_0[333] = 10'b0000001000;
assign label_0[334] = 10'b0000000010;
assign label_0[335] = 10'b0000000001;
assign label_0[336] = 10'b0000001000;
assign label_0[337] = 10'b0000000100;
assign label_0[338] = 10'b1000000000;
assign label_0[339] = 10'b0100000000;
assign label_0[340] = 10'b0000001000;
assign label_0[341] = 10'b0000001000;
assign label_0[342] = 10'b0000001000;
assign label_0[343] = 10'b0000100000;
assign label_0[344] = 10'b0100000000;
assign label_0[345] = 10'b0000001000;
assign label_0[346] = 10'b0000010000;
assign label_0[347] = 10'b1000000000;
assign label_0[348] = 10'b0100000000;
assign label_0[349] = 10'b0000001000;
assign label_0[350] = 10'b0000001000;
assign label_0[351] = 10'b0100000000;
assign label_0[352] = 10'b0000100000;
assign label_0[353] = 10'b1000000000;
assign label_0[354] = 10'b0000100000;
assign label_0[355] = 10'b0000001000;
assign label_0[356] = 10'b1000000000;
assign label_0[357] = 10'b0000001000;
assign label_0[358] = 10'b0000100000;
assign label_0[359] = 10'b1000000000;
assign label_0[360] = 10'b1000000000;
assign label_0[361] = 10'b1000000000;
assign label_0[362] = 10'b0000000100;
assign label_0[363] = 10'b0000100000;
assign label_0[364] = 10'b0000010000;
assign label_0[365] = 10'b0000001000;
assign label_0[366] = 10'b0000001000;
assign label_0[367] = 10'b0100000000;
assign label_0[368] = 10'b0000000100;
assign label_0[369] = 10'b0100000000;
assign label_0[370] = 10'b0000000100;
assign label_0[371] = 10'b0100000000;
assign label_0[372] = 10'b0100000000;
assign label_0[373] = 10'b0001000000;
assign label_0[374] = 10'b1000000000;
assign label_0[375] = 10'b0000100000;
assign label_0[376] = 10'b0000100000;
assign label_0[377] = 10'b0100000000;
assign label_0[378] = 10'b0100000000;
assign label_0[379] = 10'b0010000000;
assign label_0[380] = 10'b0000001000;
assign label_0[381] = 10'b0000100000;
assign label_0[382] = 10'b0100000000;
assign label_0[383] = 10'b0100000000;
assign label_0[384] = 10'b0000001000;
assign label_0[385] = 10'b0000001000;
assign label_0[386] = 10'b0000100000;
assign label_0[387] = 10'b0000000100;
assign label_0[388] = 10'b0000001000;
assign label_0[389] = 10'b0000001000;
assign label_0[390] = 10'b0000001000;
assign label_0[391] = 10'b0000001000;
assign label_0[392] = 10'b0000100000;
assign label_0[393] = 10'b0000100000;
assign label_0[394] = 10'b0000100000;
assign label_0[395] = 10'b0000100000;
assign label_0[396] = 10'b0000100000;
assign label_0[397] = 10'b0000100000;
assign label_0[398] = 10'b0100000000;
assign label_0[399] = 10'b0000001000;
assign label_0[400] = 10'b0000001000;
assign label_0[401] = 10'b0000000100;
assign label_0[402] = 10'b0100000000;
assign label_0[403] = 10'b0000010000;
assign label_0[404] = 10'b0000000100;
assign label_0[405] = 10'b0000000100;
assign label_0[406] = 10'b0000001000;
assign label_0[407] = 10'b0000000100;
assign label_0[408] = 10'b0000000100;
assign label_0[409] = 10'b0000001000;
assign label_0[410] = 10'b0100000000;
assign label_0[411] = 10'b0000000100;
assign label_0[412] = 10'b0000001000;
assign label_0[413] = 10'b0000010000;
assign label_0[414] = 10'b0000010000;
assign label_0[415] = 10'b0000000100;
assign label_0[416] = 10'b0000100000;
assign label_0[417] = 10'b0000100000;
assign label_0[418] = 10'b0000100000;
assign label_0[419] = 10'b0000100000;
assign label_0[420] = 10'b0000100000;
assign label_0[421] = 10'b0000100000;
assign label_0[422] = 10'b0000000100;
assign label_0[423] = 10'b0100000000;
assign label_0[424] = 10'b0000010000;
assign label_0[425] = 10'b0000010000;
assign label_0[426] = 10'b0000100000;
assign label_0[427] = 10'b1000000000;
assign label_0[428] = 10'b1000000000;
assign label_0[429] = 10'b0100000000;
assign label_0[430] = 10'b0100000000;
assign label_0[431] = 10'b1000000000;
assign label_0[432] = 10'b0000001000;
assign label_0[433] = 10'b0000001000;
assign label_0[434] = 10'b0000001000;
assign label_0[435] = 10'b0000001000;
assign label_0[436] = 10'b0000001000;
assign label_0[437] = 10'b0000001000;
assign label_0[438] = 10'b0000001000;
assign label_0[439] = 10'b0000001000;
assign label_0[440] = 10'b0000100000;
assign label_0[441] = 10'b0000100000;
assign label_0[442] = 10'b0100000000;
assign label_0[443] = 10'b0100000000;
assign label_0[444] = 10'b0000100000;
assign label_0[445] = 10'b0000100000;
assign label_0[446] = 10'b0000000001;
assign label_0[447] = 10'b0000000001;
assign label_0[448] = 10'b0000100000;
assign label_0[449] = 10'b0000100000;
assign label_0[450] = 10'b0000000001;
assign label_0[451] = 10'b0100000000;
assign label_0[452] = 10'b0000001000;
assign label_0[453] = 10'b0000001000;
assign label_0[454] = 10'b0000100000;
assign label_0[455] = 10'b0000100000;
assign label_0[456] = 10'b0000001000;
assign label_0[457] = 10'b0000100000;
assign label_0[458] = 10'b0000100000;
assign label_0[459] = 10'b0000001000;
assign label_0[460] = 10'b0000001000;
assign label_0[461] = 10'b0000001000;
assign label_0[462] = 10'b0000100000;
assign label_0[463] = 10'b0000000001;
assign label_0[464] = 10'b0000100000;
assign label_0[465] = 10'b0000001000;
assign label_0[466] = 10'b0000100000;
assign label_0[467] = 10'b0000100000;
assign label_0[468] = 10'b0000000001;
assign label_0[469] = 10'b0000000001;
assign label_0[470] = 10'b0100000000;
assign label_0[471] = 10'b0100000000;
assign label_0[472] = 10'b0000010000;
assign label_0[473] = 10'b0100000000;
assign label_0[474] = 10'b0000000001;
assign label_0[475] = 10'b0000100000;
assign label_0[476] = 10'b0000001000;
assign label_0[477] = 10'b0100000000;
assign label_0[478] = 10'b0000010000;
assign label_0[479] = 10'b0000100000;
assign label_0[480] = 10'b0000100000;
assign label_0[481] = 10'b1000000000;
assign label_0[482] = 10'b0000010000;
assign label_0[483] = 10'b0000100000;
assign label_0[484] = 10'b1000000000;
assign label_0[485] = 10'b0100000000;
assign label_0[486] = 10'b1000000000;
assign label_0[487] = 10'b0000001000;
assign label_0[488] = 10'b0000000001;
assign label_0[489] = 10'b0000100000;
assign label_0[490] = 10'b0100000000;
assign label_0[491] = 10'b1000000000;
assign label_0[492] = 10'b0000001000;
assign label_0[493] = 10'b0000001000;
assign label_0[494] = 10'b0000001000;
assign label_0[495] = 10'b0000100000;
assign label_0[496] = 10'b0100000000;
assign label_0[497] = 10'b0000000001;
assign label_0[498] = 10'b0000100000;
assign label_0[499] = 10'b0100000000;
assign label_0[500] = 10'b0000001000;
assign label_0[501] = 10'b0000100000;
assign label_0[502] = 10'b0100000000;
assign label_0[503] = 10'b0100000000;
assign label_0[504] = 10'b0000000001;
assign label_0[505] = 10'b0000000001;
assign label_0[506] = 10'b0000000100;
assign label_0[507] = 10'b0000001000;
assign label_0[508] = 10'b0100000000;
assign label_0[509] = 10'b0000001000;
assign label_0[510] = 10'b0000100000;
assign label_0[511] = 10'b0000000100;
assign label_0[512] = 10'b0000100000;
assign label_0[513] = 10'b0000000100;
assign label_0[514] = 10'b0001000000;
assign label_0[515] = 10'b0000000001;
assign label_0[516] = 10'b0000000100;
assign label_0[517] = 10'b0000000100;
assign label_0[518] = 10'b0000000001;
assign label_0[519] = 10'b0000010000;
assign label_0[520] = 10'b0000100000;
assign label_0[521] = 10'b0100000000;
assign label_0[522] = 10'b0000000100;
assign label_0[523] = 10'b0000000100;
assign label_0[524] = 10'b0000000100;
assign label_0[525] = 10'b0000000100;
assign label_0[526] = 10'b0001000000;
assign label_0[527] = 10'b0001000000;
assign label_0[528] = 10'b0001000000;
assign label_0[529] = 10'b0100000000;
assign label_0[530] = 10'b0000100000;
assign label_0[531] = 10'b0000100000;
assign label_0[532] = 10'b0000100000;
assign label_0[533] = 10'b0000100000;
assign label_0[534] = 10'b0000100000;
assign label_0[535] = 10'b0000001000;
assign label_0[536] = 10'b0000000100;
assign label_0[537] = 10'b0000001000;
assign label_0[538] = 10'b0000100000;
assign label_0[539] = 10'b0000100000;
assign label_0[540] = 10'b0100000000;
assign label_0[541] = 10'b0100000000;
assign label_0[542] = 10'b0000000010;
assign label_0[543] = 10'b0000000010;
assign label_0[544] = 10'b0000000001;
assign label_0[545] = 10'b0000000001;
assign label_0[546] = 10'b0000100000;
assign label_0[547] = 10'b0000001000;
assign label_0[548] = 10'b0000001000;
assign label_0[549] = 10'b0000000100;
assign label_0[550] = 10'b0000100000;
assign label_0[551] = 10'b0000001000;
assign label_0[552] = 10'b0000000001;
assign label_0[553] = 10'b0000000001;
assign label_0[554] = 10'b0001000000;
assign label_0[555] = 10'b0001000000;
assign label_0[556] = 10'b1000000000;
assign label_0[557] = 10'b1000000000;
assign label_0[558] = 10'b0000000001;
assign label_0[559] = 10'b0000000001;
assign label_0[560] = 10'b1000000000;
assign label_0[561] = 10'b0000000001;
assign label_0[562] = 10'b0000001000;
assign label_0[563] = 10'b0000000001;
assign label_0[564] = 10'b0000000001;
assign label_0[565] = 10'b0000000001;
assign label_0[566] = 10'b0000000001;
assign label_0[567] = 10'b0000000001;
assign label_0[568] = 10'b0000000001;
assign label_0[569] = 10'b0000000001;
assign label_0[570] = 10'b0001000000;
assign label_0[571] = 10'b0001000000;
assign label_0[572] = 10'b0001000000;
assign label_0[573] = 10'b0001000000;
assign label_0[574] = 10'b0001000000;
assign label_0[575] = 10'b0001000000;
assign label_0[576] = 10'b0001000000;
assign label_0[577] = 10'b0000000100;
assign label_0[578] = 10'b0000000010;
assign label_0[579] = 10'b0000100000;
assign label_0[580] = 10'b0000000001;
assign label_0[581] = 10'b0100000000;
assign label_0[582] = 10'b0000000100;
assign label_0[583] = 10'b0100000000;
assign label_0[584] = 10'b0000001000;
assign label_0[585] = 10'b0000000100;
assign label_0[586] = 10'b0000000100;
assign label_0[587] = 10'b0000000100;
assign label_0[588] = 10'b0100000000;
assign label_0[589] = 10'b0000001000;
assign label_0[590] = 10'b0001000000;
assign label_0[591] = 10'b0000000100;
assign label_0[592] = 10'b0000000010;
assign label_0[593] = 10'b0000000010;
assign label_0[594] = 10'b0100000000;
assign label_0[595] = 10'b0000000010;
assign label_0[596] = 10'b0000001000;
assign label_0[597] = 10'b0000000100;
assign label_0[598] = 10'b0000000100;
assign label_0[599] = 10'b0000000100;
assign label_0[600] = 10'b0000000001;
assign label_0[601] = 10'b0100000000;
assign label_0[602] = 10'b0000000100;
assign label_0[603] = 10'b0000000100;
assign label_0[604] = 10'b0100000000;
assign label_0[605] = 10'b0100000000;
assign label_0[606] = 10'b0100000000;
assign label_0[607] = 10'b0000001000;
assign label_0[608] = 10'b0000000100;
assign label_0[609] = 10'b0000000100;
assign label_0[610] = 10'b0001000000;
assign label_0[611] = 10'b0000000100;
assign label_0[612] = 10'b0010000000;
assign label_0[613] = 10'b0000000100;
assign label_0[614] = 10'b0000000001;
assign label_0[615] = 10'b0000001000;
assign label_0[616] = 10'b0100000000;
assign label_0[617] = 10'b0100000000;
assign label_0[618] = 10'b0001000000;
assign label_0[619] = 10'b0000000001;
assign label_0[620] = 10'b0000000100;
assign label_0[621] = 10'b0000000100;
assign label_0[622] = 10'b0000000100;
assign label_0[623] = 10'b0100000000;
assign label_0[624] = 10'b0000000100;
assign label_0[625] = 10'b0000000100;
assign label_0[626] = 10'b0000000100;
assign label_0[627] = 10'b0000001000;
assign label_0[628] = 10'b0000000001;
assign label_0[629] = 10'b0000000100;
assign label_0[630] = 10'b0000000100;
assign label_0[631] = 10'b0001000000;
assign label_0[632] = 10'b0001000000;
assign label_0[633] = 10'b0000000001;
assign label_0[634] = 10'b0000000100;
assign label_0[635] = 10'b0100000000;
assign label_0[636] = 10'b0000000100;
assign label_0[637] = 10'b0000000001;
assign label_0[638] = 10'b0000000100;
assign label_0[639] = 10'b0000000100;
assign label_0[640] = 10'b0001000000;
assign label_0[641] = 10'b0000010000;
assign label_0[642] = 10'b0000000001;
assign label_0[643] = 10'b0001000000;
assign label_0[644] = 10'b0000000001;
assign label_0[645] = 10'b0000000001;
assign label_0[646] = 10'b0000000001;
assign label_0[647] = 10'b0000000001;
assign label_0[648] = 10'b0000000001;
assign label_0[649] = 10'b0001000000;
assign label_0[650] = 10'b0000000100;
assign label_0[651] = 10'b0001000000;
assign label_0[652] = 10'b0000000001;
assign label_0[653] = 10'b0000000001;
assign label_0[654] = 10'b0000000100;
assign label_0[655] = 10'b0000100000;
assign label_0[656] = 10'b0010000000;
assign label_0[657] = 10'b0000000001;
assign label_0[658] = 10'b0000000001;
assign label_0[659] = 10'b0001000000;
assign label_0[660] = 10'b0001000000;
assign label_0[661] = 10'b0000000001;
assign label_0[662] = 10'b0000000001;
assign label_0[663] = 10'b0000010000;
assign label_0[664] = 10'b0000000001;
assign label_0[665] = 10'b0000000001;
assign label_0[666] = 10'b0000000001;
assign label_0[667] = 10'b0100000000;
assign label_0[668] = 10'b0000000100;
assign label_0[669] = 10'b0000000100;
assign label_0[670] = 10'b0000100000;
assign label_0[671] = 10'b0000100000;
assign label_0[672] = 10'b0000100000;
assign label_0[673] = 10'b0000001000;
assign label_0[674] = 10'b0000000001;
assign label_0[675] = 10'b0000000100;
assign label_0[676] = 10'b0000000001;
assign label_0[677] = 10'b0000000001;
assign label_0[678] = 10'b0000001000;
assign label_0[679] = 10'b0000000001;
assign label_0[680] = 10'b0000000001;
assign label_0[681] = 10'b0000100000;
assign label_0[682] = 10'b0000001000;
assign label_0[683] = 10'b0000000100;
assign label_0[684] = 10'b0000000100;
assign label_0[685] = 10'b0000000100;
assign label_0[686] = 10'b0000000100;
assign label_0[687] = 10'b0000000001;
assign label_0[688] = 10'b0000000001;
assign label_0[689] = 10'b0000000001;
assign label_0[690] = 10'b0000100000;
assign label_0[691] = 10'b0000100000;
assign label_0[692] = 10'b0000000001;
assign label_0[693] = 10'b0000000001;
assign label_0[694] = 10'b0000000001;
assign label_0[695] = 10'b0001000000;
assign label_0[696] = 10'b0000100000;
assign label_0[697] = 10'b0001000000;
assign label_0[698] = 10'b0000000001;
assign label_0[699] = 10'b0000000001;
assign label_0[700] = 10'b0000100000;
assign label_0[701] = 10'b0000000001;
assign label_0[702] = 10'b0100000000;
assign label_0[703] = 10'b0000001000;
assign label_0[704] = 10'b0000000100;
assign label_0[705] = 10'b0000010000;
assign label_0[706] = 10'b0000000100;
assign label_0[707] = 10'b0000010000;
assign label_0[708] = 10'b0000100000;
assign label_0[709] = 10'b0000010000;
assign label_0[710] = 10'b0000010000;
assign label_0[711] = 10'b0000100000;
assign label_0[712] = 10'b0001000000;
assign label_0[713] = 10'b0000000001;
assign label_0[714] = 10'b0000100000;
assign label_0[715] = 10'b0001000000;
assign label_0[716] = 10'b0000000100;
assign label_0[717] = 10'b0001000000;
assign label_0[718] = 10'b0001000000;
assign label_0[719] = 10'b0000000100;
assign label_0[720] = 10'b0000100000;
assign label_0[721] = 10'b0000000100;
assign label_0[722] = 10'b0100000000;
assign label_0[723] = 10'b0000100000;
assign label_0[724] = 10'b0000000001;
assign label_0[725] = 10'b0000000001;
assign label_0[726] = 10'b0100000000;
assign label_0[727] = 10'b0100000000;
assign label_0[728] = 10'b0000010000;
assign label_0[729] = 10'b0001000000;
assign label_0[730] = 10'b0000000001;
assign label_0[731] = 10'b0000000100;
assign label_0[732] = 10'b0000000100;
assign label_0[733] = 10'b0000000001;
assign label_0[734] = 10'b0010000000;
assign label_0[735] = 10'b1000000000;
assign label_0[736] = 10'b0000000001;
assign label_0[737] = 10'b0001000000;
assign label_0[738] = 10'b0000000100;
assign label_0[739] = 10'b0000010000;
assign label_0[740] = 10'b0000000100;
assign label_0[741] = 10'b0000000100;
assign label_0[742] = 10'b0000000100;
assign label_0[743] = 10'b0000000100;
assign label_0[744] = 10'b0001000000;
assign label_0[745] = 10'b0000100000;
assign label_0[746] = 10'b0000001000;
assign label_0[747] = 10'b0100000000;
assign label_0[748] = 10'b0000000100;
assign label_0[749] = 10'b0000000100;
assign label_0[750] = 10'b1000000000;
assign label_0[751] = 10'b0000000001;
assign label_0[752] = 10'b0001000000;
assign label_0[753] = 10'b0001000000;
assign label_0[754] = 10'b0001000000;
assign label_0[755] = 10'b0000100000;
assign label_0[756] = 10'b0001000000;
assign label_0[757] = 10'b0000100000;
assign label_0[758] = 10'b0000000100;
assign label_0[759] = 10'b0000000100;
assign label_0[760] = 10'b0000100000;
assign label_0[761] = 10'b0100000000;
assign label_0[762] = 10'b0001000000;
assign label_0[763] = 10'b0001000000;
assign label_0[764] = 10'b0000000100;
assign label_0[765] = 10'b0100000000;
assign label_0[766] = 10'b0000000001;
assign label_0[767] = 10'b0000000001;
assign label_0[768] = 10'b0001000000;
assign label_0[769] = 10'b0000010000;
assign label_0[770] = 10'b0001000000;
assign label_0[771] = 10'b0000100000;
assign label_0[772] = 10'b0000100000;
assign label_0[773] = 10'b0000001000;
assign label_0[774] = 10'b0100000000;
assign label_0[775] = 10'b0100000000;
assign label_0[776] = 10'b0000001000;
assign label_0[777] = 10'b0000100000;
assign label_0[778] = 10'b0001000000;
assign label_0[779] = 10'b0000000100;
assign label_0[780] = 10'b0000001000;
assign label_0[781] = 10'b0000100000;
assign label_0[782] = 10'b0000001000;
assign label_0[783] = 10'b0100000000;
assign label_0[784] = 10'b0000000100;
assign label_0[785] = 10'b0100000000;
assign label_0[786] = 10'b0100000000;
assign label_0[787] = 10'b1000000000;
assign label_0[788] = 10'b0001000000;
assign label_0[789] = 10'b1000000000;
assign label_0[790] = 10'b0001000000;
assign label_0[791] = 10'b0000000100;
assign label_0[792] = 10'b0000000100;
assign label_0[793] = 10'b0000000100;
assign label_0[794] = 10'b0000010000;
assign label_0[795] = 10'b1000000000;
assign label_0[796] = 10'b0000000010;
assign label_0[797] = 10'b0001000000;
assign label_0[798] = 10'b0000100000;
assign label_0[799] = 10'b0100000000;
assign label_0[800] = 10'b0000000100;
assign label_0[801] = 10'b0001000000;
assign label_0[802] = 10'b0001000000;
assign label_0[803] = 10'b0000000100;
assign label_0[804] = 10'b0001000000;
assign label_0[805] = 10'b0001000000;
assign label_0[806] = 10'b0001000000;
assign label_0[807] = 10'b0000000100;
assign label_0[808] = 10'b0000000100;
assign label_0[809] = 10'b0000010000;
assign label_0[810] = 10'b0001000000;
assign label_0[811] = 10'b0001000000;
assign label_0[812] = 10'b0000100000;
assign label_0[813] = 10'b0000100000;
assign label_0[814] = 10'b0000001000;
assign label_0[815] = 10'b0000100000;
assign label_0[816] = 10'b0000100000;
assign label_0[817] = 10'b0000100000;
assign label_0[818] = 10'b0001000000;
assign label_0[819] = 10'b0000100000;
assign label_0[820] = 10'b0100000000;
assign label_0[821] = 10'b0000010000;
assign label_0[822] = 10'b0000000100;
assign label_0[823] = 10'b0100000000;
assign label_0[824] = 10'b0000100000;
assign label_0[825] = 10'b0000000100;
assign label_0[826] = 10'b0000000100;
assign label_0[827] = 10'b0000000100;
assign label_0[828] = 10'b0000000100;
assign label_0[829] = 10'b0000000100;
assign label_0[830] = 10'b0000010000;
assign label_0[831] = 10'b0000000001;
assign label_0[832] = 10'b0100000000;
assign label_0[833] = 10'b0100000000;
assign label_0[834] = 10'b0000000100;
assign label_0[835] = 10'b0100000000;
assign label_0[836] = 10'b0000100000;
assign label_0[837] = 10'b0000100000;
assign label_0[838] = 10'b0000100000;
assign label_0[839] = 10'b0000100000;
assign label_0[840] = 10'b0000000100;
assign label_0[841] = 10'b0000000100;
assign label_0[842] = 10'b0000000100;
assign label_0[843] = 10'b0000000100;
assign label_0[844] = 10'b0000000100;
assign label_0[845] = 10'b0000000100;
assign label_0[846] = 10'b0000000100;
assign label_0[847] = 10'b0000000100;
assign label_0[848] = 10'b0100000000;
assign label_0[849] = 10'b0100000000;
assign label_0[850] = 10'b0100000000;
assign label_0[851] = 10'b0100000000;
assign label_0[852] = 10'b0000001000;
assign label_0[853] = 10'b0000001000;
assign label_0[854] = 10'b0000001000;
assign label_0[855] = 10'b0000001000;
assign label_0[856] = 10'b1000000000;
assign label_0[857] = 10'b1000000000;
assign label_0[858] = 10'b1000000000;
assign label_0[859] = 10'b1000000000;
assign label_0[860] = 10'b0000010000;
assign label_0[861] = 10'b0000010000;
assign label_0[862] = 10'b0000100000;
assign label_0[863] = 10'b0000100000;
assign label_0[864] = 10'b0000001000;
assign label_0[865] = 10'b0000001000;
assign label_0[866] = 10'b0000100000;
assign label_0[867] = 10'b0000100000;
assign label_0[868] = 10'b0000001000;
assign label_0[869] = 10'b0000100000;
assign label_0[870] = 10'b0100000000;
assign label_0[871] = 10'b0100000000;
assign label_0[872] = 10'b0100000000;
assign label_0[873] = 10'b0100000000;
assign label_0[874] = 10'b0100000000;
assign label_0[875] = 10'b0100000000;
assign label_0[876] = 10'b0100000000;
assign label_0[877] = 10'b0100000000;
assign label_0[878] = 10'b0100000000;
assign label_0[879] = 10'b0100000000;
assign label_0[880] = 10'b0000001000;
assign label_0[881] = 10'b0000100000;
assign label_0[882] = 10'b0000000100;
assign label_0[883] = 10'b0100000000;
assign label_0[884] = 10'b0100000000;
assign label_0[885] = 10'b0100000000;
assign label_0[886] = 10'b0100000000;
assign label_0[887] = 10'b0100000000;
assign label_0[888] = 10'b0000010000;
assign label_0[889] = 10'b0000010000;
assign label_0[890] = 10'b0000010000;
assign label_0[891] = 10'b0000010000;
assign label_0[892] = 10'b1000000000;
assign label_0[893] = 10'b0100000000;
assign label_0[894] = 10'b0000001000;
assign label_0[895] = 10'b0100000000;
assign label_0[896] = 10'b0000000010;
assign label_0[897] = 10'b0000000100;
assign label_0[898] = 10'b1000000000;
assign label_0[899] = 10'b0000010000;
assign label_0[900] = 10'b0000100000;
assign label_0[901] = 10'b0100000000;
assign label_0[902] = 10'b0000010000;
assign label_0[903] = 10'b0001000000;
assign label_0[904] = 10'b0000100000;
assign label_0[905] = 10'b0010000000;
assign label_0[906] = 10'b0000000010;
assign label_0[907] = 10'b0000000010;
assign label_0[908] = 10'b0010000000;
assign label_0[909] = 10'b0000100000;
assign label_0[910] = 10'b0000100000;
assign label_0[911] = 10'b0100000000;
assign label_0[912] = 10'b0000000100;
assign label_0[913] = 10'b0100000000;
assign label_0[914] = 10'b0100000000;
assign label_0[915] = 10'b1000000000;
assign label_0[916] = 10'b0000000100;
assign label_0[917] = 10'b0000000100;
assign label_0[918] = 10'b0000000100;
assign label_0[919] = 10'b0100000000;
assign label_0[920] = 10'b0000000100;
assign label_0[921] = 10'b0100000000;
assign label_0[922] = 10'b1000000000;
assign label_0[923] = 10'b0100000000;
assign label_0[924] = 10'b0100000000;
assign label_0[925] = 10'b0100000000;
assign label_0[926] = 10'b0100000000;
assign label_0[927] = 10'b0100000000;
assign label_0[928] = 10'b0000010000;
assign label_0[929] = 10'b0000100000;
assign label_0[930] = 10'b0001000000;
assign label_0[931] = 10'b0000100000;
assign label_0[932] = 10'b0000010000;
assign label_0[933] = 10'b0000000100;
assign label_0[934] = 10'b0001000000;
assign label_0[935] = 10'b0000010000;
assign label_0[936] = 10'b0000010000;
assign label_0[937] = 10'b0001000000;
assign label_0[938] = 10'b0000010000;
assign label_0[939] = 10'b0000010000;
assign label_0[940] = 10'b0001000000;
assign label_0[941] = 10'b0001000000;
assign label_0[942] = 10'b0000000001;
assign label_0[943] = 10'b0001000000;
assign label_0[944] = 10'b1000000000;
assign label_0[945] = 10'b0100000000;
assign label_0[946] = 10'b0000000100;
assign label_0[947] = 10'b0000001000;
assign label_0[948] = 10'b0000001000;
assign label_0[949] = 10'b0000000100;
assign label_0[950] = 10'b0000001000;
assign label_0[951] = 10'b0100000000;
assign label_0[952] = 10'b0000000100;
assign label_0[953] = 10'b0000000001;
assign label_0[954] = 10'b0000000100;
assign label_0[955] = 10'b0100000000;
assign label_0[956] = 10'b1000000000;
assign label_0[957] = 10'b0000010000;
assign label_0[958] = 10'b0100000000;
assign label_0[959] = 10'b0100000000;
assign label_0[960] = 10'b0000000100;
assign label_0[961] = 10'b0000000100;
assign label_0[962] = 10'b0000001000;
assign label_0[963] = 10'b0000000100;
assign label_0[964] = 10'b0000000100;
assign label_0[965] = 10'b0000000100;
assign label_0[966] = 10'b0100000000;
assign label_0[967] = 10'b0000001000;
assign label_0[968] = 10'b0000000001;
assign label_0[969] = 10'b0000000100;
assign label_0[970] = 10'b0100000000;
assign label_0[971] = 10'b0000000100;
assign label_0[972] = 10'b0000000100;
assign label_0[973] = 10'b0000000100;
assign label_0[974] = 10'b0000000001;
assign label_0[975] = 10'b0001000000;
assign label_0[976] = 10'b0000000100;
assign label_0[977] = 10'b0000000100;
assign label_0[978] = 10'b0000000100;
assign label_0[979] = 10'b0000000100;
assign label_0[980] = 10'b0000000100;
assign label_0[981] = 10'b0100000000;
assign label_0[982] = 10'b0000000100;
assign label_0[983] = 10'b0000000001;
assign label_0[984] = 10'b0100000000;
assign label_0[985] = 10'b0000000100;
assign label_0[986] = 10'b0100000000;
assign label_0[987] = 10'b0100000000;
assign label_0[988] = 10'b0000000100;
assign label_0[989] = 10'b0000000100;
assign label_0[990] = 10'b0100000000;
assign label_0[991] = 10'b0100000000;
assign label_0[992] = 10'b0000001000;
assign label_0[993] = 10'b0000001000;
assign label_0[994] = 10'b0100000000;
assign label_0[995] = 10'b0100000000;
assign label_0[996] = 10'b0100000000;
assign label_0[997] = 10'b0100000000;
assign label_0[998] = 10'b0000000001;
assign label_0[999] = 10'b0100000000;
assign label_0[1000] = 10'b0000000100;
assign label_0[1001] = 10'b0000100000;
assign label_0[1002] = 10'b0000001000;
assign label_0[1003] = 10'b0000001000;
assign label_0[1004] = 10'b0000000100;
assign label_0[1005] = 10'b0100000000;
assign label_0[1006] = 10'b0000001000;
assign label_0[1007] = 10'b0100000000;
assign label_0[1008] = 10'b0000001000;
assign label_0[1009] = 10'b0000000010;
assign label_0[1010] = 10'b0000000100;
assign label_0[1011] = 10'b0000000001;
assign label_0[1012] = 10'b0000010000;
assign label_0[1013] = 10'b0000010000;
assign label_0[1014] = 10'b0000000100;
assign label_0[1015] = 10'b0001000000;
assign label_0[1016] = 10'b0100000000;
assign label_0[1017] = 10'b0000000010;
assign label_0[1018] = 10'b0000000010;
assign label_0[1019] = 10'b0100000000;
assign label_0[1020] = 10'b0000000001;
assign label_0[1021] = 10'b0100000000;
assign label_0[1022] = 10'b0000001000;
assign label_0[1023] = 10'b0000000001;
assign label_1[0] = 10'b0000010000;
assign label_1[1] = 10'b0001000000;
assign label_1[2] = 10'b1000000000;
assign label_1[3] = 10'b0100000000;
assign label_1[4] = 10'b0000000001;
assign label_1[5] = 10'b0000000100;
assign label_1[6] = 10'b0000000100;
assign label_1[7] = 10'b0001000000;
assign label_1[8] = 10'b0000010000;
assign label_1[9] = 10'b0001000000;
assign label_1[10] = 10'b0000000001;
assign label_1[11] = 10'b0001000000;
assign label_1[12] = 10'b0001000000;
assign label_1[13] = 10'b0001000000;
assign label_1[14] = 10'b0000000001;
assign label_1[15] = 10'b0000000100;
assign label_1[16] = 10'b0000010000;
assign label_1[17] = 10'b0001000000;
assign label_1[18] = 10'b0000100000;
assign label_1[19] = 10'b0010000000;
assign label_1[20] = 10'b0000100000;
assign label_1[21] = 10'b0000100000;
assign label_1[22] = 10'b0000100000;
assign label_1[23] = 10'b0000100000;
assign label_1[24] = 10'b0000000100;
assign label_1[25] = 10'b0001000000;
assign label_1[26] = 10'b0000001000;
assign label_1[27] = 10'b0000100000;
assign label_1[28] = 10'b0000100000;
assign label_1[29] = 10'b0000100000;
assign label_1[30] = 10'b0000000001;
assign label_1[31] = 10'b0000100000;
assign label_1[32] = 10'b0000000010;
assign label_1[33] = 10'b0000000100;
assign label_1[34] = 10'b0000000100;
assign label_1[35] = 10'b0000100000;
assign label_1[36] = 10'b0010000000;
assign label_1[37] = 10'b0100000000;
assign label_1[38] = 10'b0000000100;
assign label_1[39] = 10'b0100000000;
assign label_1[40] = 10'b0000010000;
assign label_1[41] = 10'b0000000100;
assign label_1[42] = 10'b0100000000;
assign label_1[43] = 10'b1000000000;
assign label_1[44] = 10'b0001000000;
assign label_1[45] = 10'b0001000000;
assign label_1[46] = 10'b0001000000;
assign label_1[47] = 10'b0001000000;
assign label_1[48] = 10'b0000010000;
assign label_1[49] = 10'b0000000100;
assign label_1[50] = 10'b1000000000;
assign label_1[51] = 10'b0000010000;
assign label_1[52] = 10'b0001000000;
assign label_1[53] = 10'b0001000000;
assign label_1[54] = 10'b0010000000;
assign label_1[55] = 10'b0010000000;
assign label_1[56] = 10'b0010000000;
assign label_1[57] = 10'b0001000000;
assign label_1[58] = 10'b0000010000;
assign label_1[59] = 10'b0000010000;
assign label_1[60] = 10'b0001000000;
assign label_1[61] = 10'b0001000000;
assign label_1[62] = 10'b0001000000;
assign label_1[63] = 10'b0001000000;
assign label_1[64] = 10'b0000010000;
assign label_1[65] = 10'b0001000000;
assign label_1[66] = 10'b0000010000;
assign label_1[67] = 10'b0000010000;
assign label_1[68] = 10'b0001000000;
assign label_1[69] = 10'b0000010000;
assign label_1[70] = 10'b0010000000;
assign label_1[71] = 10'b1000000000;
assign label_1[72] = 10'b0000010000;
assign label_1[73] = 10'b0001000000;
assign label_1[74] = 10'b0001000000;
assign label_1[75] = 10'b0000010000;
assign label_1[76] = 10'b0000010000;
assign label_1[77] = 10'b1000000000;
assign label_1[78] = 10'b0000010000;
assign label_1[79] = 10'b1000000000;
assign label_1[80] = 10'b0001000000;
assign label_1[81] = 10'b0000010000;
assign label_1[82] = 10'b0000010000;
assign label_1[83] = 10'b0000000100;
assign label_1[84] = 10'b0001000000;
assign label_1[85] = 10'b0001000000;
assign label_1[86] = 10'b0000010000;
assign label_1[87] = 10'b0000000001;
assign label_1[88] = 10'b0000010000;
assign label_1[89] = 10'b0000000100;
assign label_1[90] = 10'b0100000000;
assign label_1[91] = 10'b0000010000;
assign label_1[92] = 10'b0000000100;
assign label_1[93] = 10'b0000000100;
assign label_1[94] = 10'b0000000001;
assign label_1[95] = 10'b0000000001;
assign label_1[96] = 10'b0000000001;
assign label_1[97] = 10'b0000010000;
assign label_1[98] = 10'b0000000100;
assign label_1[99] = 10'b0000000100;
assign label_1[100] = 10'b0000010000;
assign label_1[101] = 10'b0000010000;
assign label_1[102] = 10'b0001000000;
assign label_1[103] = 10'b0000000100;
assign label_1[104] = 10'b0100000000;
assign label_1[105] = 10'b0010000000;
assign label_1[106] = 10'b1000000000;
assign label_1[107] = 10'b0000010000;
assign label_1[108] = 10'b0000010000;
assign label_1[109] = 10'b0000010000;
assign label_1[110] = 10'b0000010000;
assign label_1[111] = 10'b0000010000;
assign label_1[112] = 10'b0000100000;
assign label_1[113] = 10'b0000010000;
assign label_1[114] = 10'b0010000000;
assign label_1[115] = 10'b0000100000;
assign label_1[116] = 10'b0010000000;
assign label_1[117] = 10'b0000010000;
assign label_1[118] = 10'b0000000100;
assign label_1[119] = 10'b0000001000;
assign label_1[120] = 10'b0000001000;
assign label_1[121] = 10'b0000001000;
assign label_1[122] = 10'b0000001000;
assign label_1[123] = 10'b0000001000;
assign label_1[124] = 10'b0000100000;
assign label_1[125] = 10'b0000010000;
assign label_1[126] = 10'b0000010000;
assign label_1[127] = 10'b0000010000;
assign label_1[128] = 10'b0010000000;
assign label_1[129] = 10'b0010000000;
assign label_1[130] = 10'b0010000000;
assign label_1[131] = 10'b0000000100;
assign label_1[132] = 10'b1000000000;
assign label_1[133] = 10'b0000000001;
assign label_1[134] = 10'b0000010000;
assign label_1[135] = 10'b0000000001;
assign label_1[136] = 10'b1000000000;
assign label_1[137] = 10'b1000000000;
assign label_1[138] = 10'b0000100000;
assign label_1[139] = 10'b0001000000;
assign label_1[140] = 10'b1000000000;
assign label_1[141] = 10'b0001000000;
assign label_1[142] = 10'b0010000000;
assign label_1[143] = 10'b1000000000;
assign label_1[144] = 10'b0010000000;
assign label_1[145] = 10'b0000010000;
assign label_1[146] = 10'b0010000000;
assign label_1[147] = 10'b0010000000;
assign label_1[148] = 10'b0010000000;
assign label_1[149] = 10'b0000100000;
assign label_1[150] = 10'b1000000000;
assign label_1[151] = 10'b0010000000;
assign label_1[152] = 10'b0000100000;
assign label_1[153] = 10'b1000000000;
assign label_1[154] = 10'b0000010000;
assign label_1[155] = 10'b1000000000;
assign label_1[156] = 10'b1000000000;
assign label_1[157] = 10'b0000010000;
assign label_1[158] = 10'b0000010000;
assign label_1[159] = 10'b1000000000;
assign label_1[160] = 10'b0001000000;
assign label_1[161] = 10'b0000000100;
assign label_1[162] = 10'b0000000001;
assign label_1[163] = 10'b0000100000;
assign label_1[164] = 10'b0000000001;
assign label_1[165] = 10'b0000000100;
assign label_1[166] = 10'b0000100000;
assign label_1[167] = 10'b0100000000;
assign label_1[168] = 10'b0000000001;
assign label_1[169] = 10'b0000000100;
assign label_1[170] = 10'b0100000000;
assign label_1[171] = 10'b0000000100;
assign label_1[172] = 10'b0000000100;
assign label_1[173] = 10'b0010000000;
assign label_1[174] = 10'b0100000000;
assign label_1[175] = 10'b0001000000;
assign label_1[176] = 10'b0000100000;
assign label_1[177] = 10'b0000000100;
assign label_1[178] = 10'b0000100000;
assign label_1[179] = 10'b0001000000;
assign label_1[180] = 10'b0010000000;
assign label_1[181] = 10'b0100000000;
assign label_1[182] = 10'b0010000000;
assign label_1[183] = 10'b0100000000;
assign label_1[184] = 10'b0000100000;
assign label_1[185] = 10'b0000000001;
assign label_1[186] = 10'b0000010000;
assign label_1[187] = 10'b0100000000;
assign label_1[188] = 10'b0000000001;
assign label_1[189] = 10'b0001000000;
assign label_1[190] = 10'b0000000001;
assign label_1[191] = 10'b0001000000;
assign label_1[192] = 10'b0000000100;
assign label_1[193] = 10'b1000000000;
assign label_1[194] = 10'b0000000001;
assign label_1[195] = 10'b0000000100;
assign label_1[196] = 10'b0000100000;
assign label_1[197] = 10'b0000100000;
assign label_1[198] = 10'b0000000001;
assign label_1[199] = 10'b0001000000;
assign label_1[200] = 10'b0000000001;
assign label_1[201] = 10'b0000000001;
assign label_1[202] = 10'b0010000000;
assign label_1[203] = 10'b0010000000;
assign label_1[204] = 10'b1000000000;
assign label_1[205] = 10'b0000000001;
assign label_1[206] = 10'b0010000000;
assign label_1[207] = 10'b1000000000;
assign label_1[208] = 10'b1000000000;
assign label_1[209] = 10'b0000000100;
assign label_1[210] = 10'b0000010000;
assign label_1[211] = 10'b0001000000;
assign label_1[212] = 10'b0000000100;
assign label_1[213] = 10'b1000000000;
assign label_1[214] = 10'b0000010000;
assign label_1[215] = 10'b1000000000;
assign label_1[216] = 10'b0000010000;
assign label_1[217] = 10'b0000000100;
assign label_1[218] = 10'b0000010000;
assign label_1[219] = 10'b0001000000;
assign label_1[220] = 10'b1000000000;
assign label_1[221] = 10'b0001000000;
assign label_1[222] = 10'b0000000100;
assign label_1[223] = 10'b1000000000;
assign label_1[224] = 10'b0000000001;
assign label_1[225] = 10'b0000000001;
assign label_1[226] = 10'b0001000000;
assign label_1[227] = 10'b0000000001;
assign label_1[228] = 10'b0100000000;
assign label_1[229] = 10'b0000000100;
assign label_1[230] = 10'b0000000001;
assign label_1[231] = 10'b0000010000;
assign label_1[232] = 10'b0000100000;
assign label_1[233] = 10'b0001000000;
assign label_1[234] = 10'b0000000001;
assign label_1[235] = 10'b0000000100;
assign label_1[236] = 10'b0000000001;
assign label_1[237] = 10'b0001000000;
assign label_1[238] = 10'b0000000100;
assign label_1[239] = 10'b0000000001;
assign label_1[240] = 10'b0000000100;
assign label_1[241] = 10'b0010000000;
assign label_1[242] = 10'b0000000100;
assign label_1[243] = 10'b0100000000;
assign label_1[244] = 10'b0000000100;
assign label_1[245] = 10'b0000000100;
assign label_1[246] = 10'b0000000100;
assign label_1[247] = 10'b0000000001;
assign label_1[248] = 10'b0000100000;
assign label_1[249] = 10'b0000000001;
assign label_1[250] = 10'b0000000001;
assign label_1[251] = 10'b0000000001;
assign label_1[252] = 10'b0000100000;
assign label_1[253] = 10'b0001000000;
assign label_1[254] = 10'b0001000000;
assign label_1[255] = 10'b0100000000;
assign label_1[256] = 10'b0000001000;
assign label_1[257] = 10'b0000100000;
assign label_1[258] = 10'b1000000000;
assign label_1[259] = 10'b1000000000;
assign label_1[260] = 10'b0001000000;
assign label_1[261] = 10'b0000000100;
assign label_1[262] = 10'b0000000001;
assign label_1[263] = 10'b0000100000;
assign label_1[264] = 10'b0000100000;
assign label_1[265] = 10'b0000000001;
assign label_1[266] = 10'b0000000001;
assign label_1[267] = 10'b0000000100;
assign label_1[268] = 10'b0000000001;
assign label_1[269] = 10'b0000000001;
assign label_1[270] = 10'b0000000100;
assign label_1[271] = 10'b0000000100;
assign label_1[272] = 10'b0000000100;
assign label_1[273] = 10'b0000000100;
assign label_1[274] = 10'b0000000010;
assign label_1[275] = 10'b0000000100;
assign label_1[276] = 10'b0000000100;
assign label_1[277] = 10'b0001000000;
assign label_1[278] = 10'b0001000000;
assign label_1[279] = 10'b0000010000;
assign label_1[280] = 10'b0001000000;
assign label_1[281] = 10'b0000000100;
assign label_1[282] = 10'b0001000000;
assign label_1[283] = 10'b0000001000;
assign label_1[284] = 10'b0000010000;
assign label_1[285] = 10'b0001000000;
assign label_1[286] = 10'b0100000000;
assign label_1[287] = 10'b0000100000;
assign label_1[288] = 10'b0000000001;
assign label_1[289] = 10'b0000000001;
assign label_1[290] = 10'b0000001000;
assign label_1[291] = 10'b0000001000;
assign label_1[292] = 10'b0000000001;
assign label_1[293] = 10'b0000000001;
assign label_1[294] = 10'b0000001000;
assign label_1[295] = 10'b0000000100;
assign label_1[296] = 10'b0000000100;
assign label_1[297] = 10'b0000000001;
assign label_1[298] = 10'b0000001000;
assign label_1[299] = 10'b0000000100;
assign label_1[300] = 10'b0000000100;
assign label_1[301] = 10'b0000000001;
assign label_1[302] = 10'b0000000001;
assign label_1[303] = 10'b0000000001;
assign label_1[304] = 10'b0000000100;
assign label_1[305] = 10'b0000000100;
assign label_1[306] = 10'b0000000100;
assign label_1[307] = 10'b0000100000;
assign label_1[308] = 10'b0100000000;
assign label_1[309] = 10'b0001000000;
assign label_1[310] = 10'b0000010000;
assign label_1[311] = 10'b0000100000;
assign label_1[312] = 10'b0000010000;
assign label_1[313] = 10'b0000010000;
assign label_1[314] = 10'b1000000000;
assign label_1[315] = 10'b0000001000;
assign label_1[316] = 10'b0100000000;
assign label_1[317] = 10'b0100000000;
assign label_1[318] = 10'b0000100000;
assign label_1[319] = 10'b0000100000;
assign label_1[320] = 10'b0000000001;
assign label_1[321] = 10'b0000100000;
assign label_1[322] = 10'b0000000001;
assign label_1[323] = 10'b0001000000;
assign label_1[324] = 10'b0000000001;
assign label_1[325] = 10'b0000100000;
assign label_1[326] = 10'b0000000001;
assign label_1[327] = 10'b0000000001;
assign label_1[328] = 10'b0000000001;
assign label_1[329] = 10'b0000000001;
assign label_1[330] = 10'b0000001000;
assign label_1[331] = 10'b0000001000;
assign label_1[332] = 10'b0001000000;
assign label_1[333] = 10'b0000000100;
assign label_1[334] = 10'b0001000000;
assign label_1[335] = 10'b0000000001;
assign label_1[336] = 10'b0001000000;
assign label_1[337] = 10'b0000000001;
assign label_1[338] = 10'b0000100000;
assign label_1[339] = 10'b0000000010;
assign label_1[340] = 10'b0001000000;
assign label_1[341] = 10'b0001000000;
assign label_1[342] = 10'b0000000001;
assign label_1[343] = 10'b0000000001;
assign label_1[344] = 10'b1000000000;
assign label_1[345] = 10'b0000010000;
assign label_1[346] = 10'b0001000000;
assign label_1[347] = 10'b0000000001;
assign label_1[348] = 10'b0000001000;
assign label_1[349] = 10'b0000100000;
assign label_1[350] = 10'b0000000001;
assign label_1[351] = 10'b0000000001;
assign label_1[352] = 10'b0000100000;
assign label_1[353] = 10'b0001000000;
assign label_1[354] = 10'b0000100000;
assign label_1[355] = 10'b0000100000;
assign label_1[356] = 10'b1000000000;
assign label_1[357] = 10'b0000010000;
assign label_1[358] = 10'b0001000000;
assign label_1[359] = 10'b0000000100;
assign label_1[360] = 10'b0000000001;
assign label_1[361] = 10'b0000000001;
assign label_1[362] = 10'b0001000000;
assign label_1[363] = 10'b0001000000;
assign label_1[364] = 10'b0000010000;
assign label_1[365] = 10'b0000010000;
assign label_1[366] = 10'b0100000000;
assign label_1[367] = 10'b0000000100;
assign label_1[368] = 10'b0000100000;
assign label_1[369] = 10'b0000100000;
assign label_1[370] = 10'b0000010000;
assign label_1[371] = 10'b0000100000;
assign label_1[372] = 10'b0001000000;
assign label_1[373] = 10'b0000100000;
assign label_1[374] = 10'b0000000001;
assign label_1[375] = 10'b0000000001;
assign label_1[376] = 10'b0100000000;
assign label_1[377] = 10'b0100000000;
assign label_1[378] = 10'b0100000000;
assign label_1[379] = 10'b0100000000;
assign label_1[380] = 10'b0000000001;
assign label_1[381] = 10'b1000000000;
assign label_1[382] = 10'b1000000000;
assign label_1[383] = 10'b0000000001;
assign label_1[384] = 10'b0000010000;
assign label_1[385] = 10'b0000000100;
assign label_1[386] = 10'b1000000000;
assign label_1[387] = 10'b0100000000;
assign label_1[388] = 10'b0000010000;
assign label_1[389] = 10'b0000100000;
assign label_1[390] = 10'b0000010000;
assign label_1[391] = 10'b0000010000;
assign label_1[392] = 10'b0000010000;
assign label_1[393] = 10'b0000010000;
assign label_1[394] = 10'b1000000000;
assign label_1[395] = 10'b0000010000;
assign label_1[396] = 10'b0000001000;
assign label_1[397] = 10'b0000001000;
assign label_1[398] = 10'b0000000001;
assign label_1[399] = 10'b0000000100;
assign label_1[400] = 10'b0100000000;
assign label_1[401] = 10'b0000001000;
assign label_1[402] = 10'b0000100000;
assign label_1[403] = 10'b0000001000;
assign label_1[404] = 10'b0000001000;
assign label_1[405] = 10'b0000001000;
assign label_1[406] = 10'b0000001000;
assign label_1[407] = 10'b0000001000;
assign label_1[408] = 10'b0100000000;
assign label_1[409] = 10'b0100000000;
assign label_1[410] = 10'b0000000100;
assign label_1[411] = 10'b0100000000;
assign label_1[412] = 10'b0000100000;
assign label_1[413] = 10'b0000100000;
assign label_1[414] = 10'b0000100000;
assign label_1[415] = 10'b0000100000;
assign label_1[416] = 10'b0001000000;
assign label_1[417] = 10'b0001000000;
assign label_1[418] = 10'b0000000001;
assign label_1[419] = 10'b0000000100;
assign label_1[420] = 10'b0001000000;
assign label_1[421] = 10'b0000010000;
assign label_1[422] = 10'b0100000000;
assign label_1[423] = 10'b0100000000;
assign label_1[424] = 10'b0000000100;
assign label_1[425] = 10'b0000000100;
assign label_1[426] = 10'b0000000010;
assign label_1[427] = 10'b0000000100;
assign label_1[428] = 10'b0001000000;
assign label_1[429] = 10'b0000000100;
assign label_1[430] = 10'b0000000100;
assign label_1[431] = 10'b0001000000;
assign label_1[432] = 10'b0000000100;
assign label_1[433] = 10'b0000000100;
assign label_1[434] = 10'b0000001000;
assign label_1[435] = 10'b0000000100;
assign label_1[436] = 10'b0010000000;
assign label_1[437] = 10'b1000000000;
assign label_1[438] = 10'b0000000100;
assign label_1[439] = 10'b0100000000;
assign label_1[440] = 10'b0100000000;
assign label_1[441] = 10'b0000010000;
assign label_1[442] = 10'b0100000000;
assign label_1[443] = 10'b0000000100;
assign label_1[444] = 10'b0001000000;
assign label_1[445] = 10'b0000010000;
assign label_1[446] = 10'b0100000000;
assign label_1[447] = 10'b1000000000;
assign label_1[448] = 10'b0000000100;
assign label_1[449] = 10'b0100000000;
assign label_1[450] = 10'b0000000100;
assign label_1[451] = 10'b0000000001;
assign label_1[452] = 10'b0000000100;
assign label_1[453] = 10'b0001000000;
assign label_1[454] = 10'b0100000000;
assign label_1[455] = 10'b0000000100;
assign label_1[456] = 10'b0000000100;
assign label_1[457] = 10'b0000000100;
assign label_1[458] = 10'b0000010000;
assign label_1[459] = 10'b0001000000;
assign label_1[460] = 10'b0000000100;
assign label_1[461] = 10'b0000000001;
assign label_1[462] = 10'b0100000000;
assign label_1[463] = 10'b0100000000;
assign label_1[464] = 10'b0001000000;
assign label_1[465] = 10'b0000000001;
assign label_1[466] = 10'b0000000001;
assign label_1[467] = 10'b0000100000;
assign label_1[468] = 10'b0000001000;
assign label_1[469] = 10'b0000001000;
assign label_1[470] = 10'b0000001000;
assign label_1[471] = 10'b0000000100;
assign label_1[472] = 10'b0000000100;
assign label_1[473] = 10'b0000000100;
assign label_1[474] = 10'b0100000000;
assign label_1[475] = 10'b0100000000;
assign label_1[476] = 10'b0000001000;
assign label_1[477] = 10'b0000001000;
assign label_1[478] = 10'b0100000000;
assign label_1[479] = 10'b0000010000;
assign label_1[480] = 10'b0001000000;
assign label_1[481] = 10'b0000100000;
assign label_1[482] = 10'b0001000000;
assign label_1[483] = 10'b0000000100;
assign label_1[484] = 10'b0000000100;
assign label_1[485] = 10'b0000000100;
assign label_1[486] = 10'b0000000001;
assign label_1[487] = 10'b0000001000;
assign label_1[488] = 10'b0000100000;
assign label_1[489] = 10'b0100000000;
assign label_1[490] = 10'b0000100000;
assign label_1[491] = 10'b0000000100;
assign label_1[492] = 10'b0000001000;
assign label_1[493] = 10'b0000000100;
assign label_1[494] = 10'b0000000001;
assign label_1[495] = 10'b0100000000;
assign label_1[496] = 10'b0000000100;
assign label_1[497] = 10'b0000000100;
assign label_1[498] = 10'b0000000100;
assign label_1[499] = 10'b0001000000;
assign label_1[500] = 10'b0000000100;
assign label_1[501] = 10'b0001000000;
assign label_1[502] = 10'b0100000000;
assign label_1[503] = 10'b0000000001;
assign label_1[504] = 10'b0000000001;
assign label_1[505] = 10'b0000000100;
assign label_1[506] = 10'b0000000001;
assign label_1[507] = 10'b0000000100;
assign label_1[508] = 10'b0000000100;
assign label_1[509] = 10'b0000000100;
assign label_1[510] = 10'b0000000001;
assign label_1[511] = 10'b0100000000;
assign label_1[512] = 10'b0000000010;
assign label_1[513] = 10'b0000100000;
assign label_1[514] = 10'b1000000000;
assign label_1[515] = 10'b0000100000;
assign label_1[516] = 10'b0000100000;
assign label_1[517] = 10'b0000001000;
assign label_1[518] = 10'b0000001000;
assign label_1[519] = 10'b0001000000;
assign label_1[520] = 10'b0000100000;
assign label_1[521] = 10'b0000100000;
assign label_1[522] = 10'b0000100000;
assign label_1[523] = 10'b0000001000;
assign label_1[524] = 10'b0000001000;
assign label_1[525] = 10'b0000001000;
assign label_1[526] = 10'b0100000000;
assign label_1[527] = 10'b0100000000;
assign label_1[528] = 10'b0010000000;
assign label_1[529] = 10'b0000100000;
assign label_1[530] = 10'b1000000000;
assign label_1[531] = 10'b0000100000;
assign label_1[532] = 10'b0100000000;
assign label_1[533] = 10'b1000000000;
assign label_1[534] = 10'b0000001000;
assign label_1[535] = 10'b0000001000;
assign label_1[536] = 10'b0000001000;
assign label_1[537] = 10'b0100000000;
assign label_1[538] = 10'b0100000000;
assign label_1[539] = 10'b0000100000;
assign label_1[540] = 10'b0000001000;
assign label_1[541] = 10'b0000001000;
assign label_1[542] = 10'b0000001000;
assign label_1[543] = 10'b0000001000;
assign label_1[544] = 10'b1000000000;
assign label_1[545] = 10'b0000000001;
assign label_1[546] = 10'b0000100000;
assign label_1[547] = 10'b0000000100;
assign label_1[548] = 10'b0000000001;
assign label_1[549] = 10'b0000000001;
assign label_1[550] = 10'b0000000100;
assign label_1[551] = 10'b0000000001;
assign label_1[552] = 10'b0000100000;
assign label_1[553] = 10'b0000100000;
assign label_1[554] = 10'b1000000000;
assign label_1[555] = 10'b1000000000;
assign label_1[556] = 10'b0000001000;
assign label_1[557] = 10'b0000100000;
assign label_1[558] = 10'b0000100000;
assign label_1[559] = 10'b0000000001;
assign label_1[560] = 10'b0000100000;
assign label_1[561] = 10'b0000001000;
assign label_1[562] = 10'b1000000000;
assign label_1[563] = 10'b0000010000;
assign label_1[564] = 10'b0000000001;
assign label_1[565] = 10'b0000000001;
assign label_1[566] = 10'b0010000000;
assign label_1[567] = 10'b0000000001;
assign label_1[568] = 10'b1000000000;
assign label_1[569] = 10'b0000000001;
assign label_1[570] = 10'b0010000000;
assign label_1[571] = 10'b0000000001;
assign label_1[572] = 10'b0010000000;
assign label_1[573] = 10'b0000001000;
assign label_1[574] = 10'b0010000000;
assign label_1[575] = 10'b0100000000;
assign label_1[576] = 10'b0000000010;
assign label_1[577] = 10'b0000000100;
assign label_1[578] = 10'b0000000010;
assign label_1[579] = 10'b0100000000;
assign label_1[580] = 10'b0000000010;
assign label_1[581] = 10'b0000010000;
assign label_1[582] = 10'b1000000000;
assign label_1[583] = 10'b0000000100;
assign label_1[584] = 10'b0000000010;
assign label_1[585] = 10'b0000000100;
assign label_1[586] = 10'b0000000100;
assign label_1[587] = 10'b1000000000;
assign label_1[588] = 10'b0000001000;
assign label_1[589] = 10'b0000000100;
assign label_1[590] = 10'b0100000000;
assign label_1[591] = 10'b0100000000;
assign label_1[592] = 10'b0000000010;
assign label_1[593] = 10'b0100000000;
assign label_1[594] = 10'b0100000000;
assign label_1[595] = 10'b0000001000;
assign label_1[596] = 10'b0001000000;
assign label_1[597] = 10'b0001000000;
assign label_1[598] = 10'b0001000000;
assign label_1[599] = 10'b0001000000;
assign label_1[600] = 10'b0000000010;
assign label_1[601] = 10'b0000000100;
assign label_1[602] = 10'b0000001000;
assign label_1[603] = 10'b0001000000;
assign label_1[604] = 10'b0001000000;
assign label_1[605] = 10'b0001000000;
assign label_1[606] = 10'b0000000001;
assign label_1[607] = 10'b0000000001;
assign label_1[608] = 10'b1000000000;
assign label_1[609] = 10'b0000001000;
assign label_1[610] = 10'b0100000000;
assign label_1[611] = 10'b0000000001;
assign label_1[612] = 10'b0000000010;
assign label_1[613] = 10'b0000100000;
assign label_1[614] = 10'b0100000000;
assign label_1[615] = 10'b0001000000;
assign label_1[616] = 10'b0000000010;
assign label_1[617] = 10'b0000000010;
assign label_1[618] = 10'b0000100000;
assign label_1[619] = 10'b0100000000;
assign label_1[620] = 10'b0000001000;
assign label_1[621] = 10'b1000000000;
assign label_1[622] = 10'b0100000000;
assign label_1[623] = 10'b0001000000;
assign label_1[624] = 10'b0000000010;
assign label_1[625] = 10'b0100000000;
assign label_1[626] = 10'b0000000100;
assign label_1[627] = 10'b0000000100;
assign label_1[628] = 10'b0100000000;
assign label_1[629] = 10'b0000000100;
assign label_1[630] = 10'b0000000100;
assign label_1[631] = 10'b0100000000;
assign label_1[632] = 10'b0100000000;
assign label_1[633] = 10'b1000000000;
assign label_1[634] = 10'b0100000000;
assign label_1[635] = 10'b0001000000;
assign label_1[636] = 10'b0001000000;
assign label_1[637] = 10'b0001000000;
assign label_1[638] = 10'b0001000000;
assign label_1[639] = 10'b0001000000;
assign label_1[640] = 10'b0000100000;
assign label_1[641] = 10'b0000010000;
assign label_1[642] = 10'b0000100000;
assign label_1[643] = 10'b0000100000;
assign label_1[644] = 10'b1000000000;
assign label_1[645] = 10'b0100000000;
assign label_1[646] = 10'b0000001000;
assign label_1[647] = 10'b0000001000;
assign label_1[648] = 10'b1000000000;
assign label_1[649] = 10'b0000010000;
assign label_1[650] = 10'b0000010000;
assign label_1[651] = 10'b0000100000;
assign label_1[652] = 10'b0000100000;
assign label_1[653] = 10'b0001000000;
assign label_1[654] = 10'b1000000000;
assign label_1[655] = 10'b0000100000;
assign label_1[656] = 10'b0000100000;
assign label_1[657] = 10'b0000001000;
assign label_1[658] = 10'b0000100000;
assign label_1[659] = 10'b0000100000;
assign label_1[660] = 10'b0000100000;
assign label_1[661] = 10'b0000000001;
assign label_1[662] = 10'b0000001000;
assign label_1[663] = 10'b0100000000;
assign label_1[664] = 10'b0000100000;
assign label_1[665] = 10'b0100000000;
assign label_1[666] = 10'b0000100000;
assign label_1[667] = 10'b0000100000;
assign label_1[668] = 10'b0100000000;
assign label_1[669] = 10'b0000000001;
assign label_1[670] = 10'b0100000000;
assign label_1[671] = 10'b0100000000;
assign label_1[672] = 10'b0000000010;
assign label_1[673] = 10'b0000000100;
assign label_1[674] = 10'b0001000000;
assign label_1[675] = 10'b0100000000;
assign label_1[676] = 10'b0000000100;
assign label_1[677] = 10'b0000000100;
assign label_1[678] = 10'b0010000000;
assign label_1[679] = 10'b0000000100;
assign label_1[680] = 10'b0001000000;
assign label_1[681] = 10'b0000100000;
assign label_1[682] = 10'b0000100000;
assign label_1[683] = 10'b0100000000;
assign label_1[684] = 10'b0000010000;
assign label_1[685] = 10'b0100000000;
assign label_1[686] = 10'b0100000000;
assign label_1[687] = 10'b0100000000;
assign label_1[688] = 10'b0000000010;
assign label_1[689] = 10'b0100000000;
assign label_1[690] = 10'b0000010000;
assign label_1[691] = 10'b0100000000;
assign label_1[692] = 10'b0000010000;
assign label_1[693] = 10'b0001000000;
assign label_1[694] = 10'b0000010000;
assign label_1[695] = 10'b0010000000;
assign label_1[696] = 10'b0100000000;
assign label_1[697] = 10'b0000001000;
assign label_1[698] = 10'b0000001000;
assign label_1[699] = 10'b0000000001;
assign label_1[700] = 10'b0100000000;
assign label_1[701] = 10'b0000000100;
assign label_1[702] = 10'b0100000000;
assign label_1[703] = 10'b0100000000;
assign label_1[704] = 10'b0000100000;
assign label_1[705] = 10'b0001000000;
assign label_1[706] = 10'b0000100000;
assign label_1[707] = 10'b0000000100;
assign label_1[708] = 10'b0000001000;
assign label_1[709] = 10'b0000000100;
assign label_1[710] = 10'b0000100000;
assign label_1[711] = 10'b0000001000;
assign label_1[712] = 10'b0000000100;
assign label_1[713] = 10'b0000000100;
assign label_1[714] = 10'b0000001000;
assign label_1[715] = 10'b0000001000;
assign label_1[716] = 10'b0000010000;
assign label_1[717] = 10'b0000010000;
assign label_1[718] = 10'b0000000100;
assign label_1[719] = 10'b0000000100;
assign label_1[720] = 10'b0100000000;
assign label_1[721] = 10'b0000001000;
assign label_1[722] = 10'b0000000100;
assign label_1[723] = 10'b0000000100;
assign label_1[724] = 10'b0000000100;
assign label_1[725] = 10'b0000000100;
assign label_1[726] = 10'b0000000100;
assign label_1[727] = 10'b0000001000;
assign label_1[728] = 10'b0000000100;
assign label_1[729] = 10'b0000000100;
assign label_1[730] = 10'b0000001000;
assign label_1[731] = 10'b0000000100;
assign label_1[732] = 10'b0000001000;
assign label_1[733] = 10'b0000001000;
assign label_1[734] = 10'b0000000100;
assign label_1[735] = 10'b0100000000;
assign label_1[736] = 10'b1000000000;
assign label_1[737] = 10'b1000000000;
assign label_1[738] = 10'b0001000000;
assign label_1[739] = 10'b0001000000;
assign label_1[740] = 10'b0001000000;
assign label_1[741] = 10'b0001000000;
assign label_1[742] = 10'b0001000000;
assign label_1[743] = 10'b0001000000;
assign label_1[744] = 10'b0000000100;
assign label_1[745] = 10'b0000000100;
assign label_1[746] = 10'b0000001000;
assign label_1[747] = 10'b0000001000;
assign label_1[748] = 10'b0001000000;
assign label_1[749] = 10'b0001000000;
assign label_1[750] = 10'b0000000001;
assign label_1[751] = 10'b0000000001;
assign label_1[752] = 10'b0001000000;
assign label_1[753] = 10'b0100000000;
assign label_1[754] = 10'b0001000000;
assign label_1[755] = 10'b0001000000;
assign label_1[756] = 10'b0001000000;
assign label_1[757] = 10'b0000000100;
assign label_1[758] = 10'b0000100000;
assign label_1[759] = 10'b0000001000;
assign label_1[760] = 10'b0000000100;
assign label_1[761] = 10'b0000000100;
assign label_1[762] = 10'b0000000100;
assign label_1[763] = 10'b0000000100;
assign label_1[764] = 10'b0000000100;
assign label_1[765] = 10'b0000000100;
assign label_1[766] = 10'b0001000000;
assign label_1[767] = 10'b0001000000;
assign label_1[768] = 10'b0000010000;
assign label_1[769] = 10'b0000001000;
assign label_1[770] = 10'b0000000100;
assign label_1[771] = 10'b0001000000;
assign label_1[772] = 10'b0000001000;
assign label_1[773] = 10'b0100000000;
assign label_1[774] = 10'b0000100000;
assign label_1[775] = 10'b0000010000;
assign label_1[776] = 10'b0000001000;
assign label_1[777] = 10'b0000001000;
assign label_1[778] = 10'b0000000001;
assign label_1[779] = 10'b0000100000;
assign label_1[780] = 10'b0000000100;
assign label_1[781] = 10'b0000010000;
assign label_1[782] = 10'b0000001000;
assign label_1[783] = 10'b0000001000;
assign label_1[784] = 10'b0000010000;
assign label_1[785] = 10'b0100000000;
assign label_1[786] = 10'b0000100000;
assign label_1[787] = 10'b0000001000;
assign label_1[788] = 10'b0000001000;
assign label_1[789] = 10'b0000100000;
assign label_1[790] = 10'b0000100000;
assign label_1[791] = 10'b0000010000;
assign label_1[792] = 10'b0001000000;
assign label_1[793] = 10'b0001000000;
assign label_1[794] = 10'b0000000100;
assign label_1[795] = 10'b0001000000;
assign label_1[796] = 10'b0000000100;
assign label_1[797] = 10'b0100000000;
assign label_1[798] = 10'b0000100000;
assign label_1[799] = 10'b0000100000;
assign label_1[800] = 10'b0000001000;
assign label_1[801] = 10'b0000000100;
assign label_1[802] = 10'b0000000100;
assign label_1[803] = 10'b0001000000;
assign label_1[804] = 10'b0000001000;
assign label_1[805] = 10'b0000000100;
assign label_1[806] = 10'b0000100000;
assign label_1[807] = 10'b0000001000;
assign label_1[808] = 10'b0000100000;
assign label_1[809] = 10'b0100000000;
assign label_1[810] = 10'b0000100000;
assign label_1[811] = 10'b1000000000;
assign label_1[812] = 10'b0000000100;
assign label_1[813] = 10'b0100000000;
assign label_1[814] = 10'b0000001000;
assign label_1[815] = 10'b0000001000;
assign label_1[816] = 10'b0000001000;
assign label_1[817] = 10'b0000100000;
assign label_1[818] = 10'b0000001000;
assign label_1[819] = 10'b0000001000;
assign label_1[820] = 10'b1000000000;
assign label_1[821] = 10'b0000001000;
assign label_1[822] = 10'b0000100000;
assign label_1[823] = 10'b0000100000;
assign label_1[824] = 10'b0000001000;
assign label_1[825] = 10'b0000001000;
assign label_1[826] = 10'b0000100000;
assign label_1[827] = 10'b0100000000;
assign label_1[828] = 10'b0000000100;
assign label_1[829] = 10'b0100000000;
assign label_1[830] = 10'b0001000000;
assign label_1[831] = 10'b0100000000;
assign label_1[832] = 10'b0000100000;
assign label_1[833] = 10'b0000100000;
assign label_1[834] = 10'b0000000010;
assign label_1[835] = 10'b0000010000;
assign label_1[836] = 10'b0000001000;
assign label_1[837] = 10'b0000100000;
assign label_1[838] = 10'b0000000100;
assign label_1[839] = 10'b0100000000;
assign label_1[840] = 10'b0000010000;
assign label_1[841] = 10'b1000000000;
assign label_1[842] = 10'b0100000000;
assign label_1[843] = 10'b0000000001;
assign label_1[844] = 10'b0000100000;
assign label_1[845] = 10'b0000000001;
assign label_1[846] = 10'b0000001000;
assign label_1[847] = 10'b0000001000;
assign label_1[848] = 10'b0001000000;
assign label_1[849] = 10'b0001000000;
assign label_1[850] = 10'b0000000001;
assign label_1[851] = 10'b0001000000;
assign label_1[852] = 10'b0100000000;
assign label_1[853] = 10'b0100000000;
assign label_1[854] = 10'b0000010000;
assign label_1[855] = 10'b0000100000;
assign label_1[856] = 10'b0100000000;
assign label_1[857] = 10'b0100000000;
assign label_1[858] = 10'b0100000000;
assign label_1[859] = 10'b0000100000;
assign label_1[860] = 10'b0000100000;
assign label_1[861] = 10'b0000001000;
assign label_1[862] = 10'b0100000000;
assign label_1[863] = 10'b0000000001;
assign label_1[864] = 10'b0100000000;
assign label_1[865] = 10'b0100000000;
assign label_1[866] = 10'b0000001000;
assign label_1[867] = 10'b0000001000;
assign label_1[868] = 10'b0000001000;
assign label_1[869] = 10'b0000001000;
assign label_1[870] = 10'b0000001000;
assign label_1[871] = 10'b0000001000;
assign label_1[872] = 10'b0000100000;
assign label_1[873] = 10'b0000001000;
assign label_1[874] = 10'b0000001000;
assign label_1[875] = 10'b0000000001;
assign label_1[876] = 10'b0000100000;
assign label_1[877] = 10'b0000010000;
assign label_1[878] = 10'b0000001000;
assign label_1[879] = 10'b0000001000;
assign label_1[880] = 10'b0000000100;
assign label_1[881] = 10'b0100000000;
assign label_1[882] = 10'b0000001000;
assign label_1[883] = 10'b0000001000;
assign label_1[884] = 10'b0000001000;
assign label_1[885] = 10'b0100000000;
assign label_1[886] = 10'b0000000100;
assign label_1[887] = 10'b0000000001;
assign label_1[888] = 10'b0000100000;
assign label_1[889] = 10'b0000100000;
assign label_1[890] = 10'b0000100000;
assign label_1[891] = 10'b0000100000;
assign label_1[892] = 10'b0000100000;
assign label_1[893] = 10'b0000100000;
assign label_1[894] = 10'b0000100000;
assign label_1[895] = 10'b0000100000;
assign label_1[896] = 10'b0000001000;
assign label_1[897] = 10'b0000000100;
assign label_1[898] = 10'b0000000010;
assign label_1[899] = 10'b0100000000;
assign label_1[900] = 10'b0000001000;
assign label_1[901] = 10'b0000001000;
assign label_1[902] = 10'b0100000000;
assign label_1[903] = 10'b0000001000;
assign label_1[904] = 10'b0000000100;
assign label_1[905] = 10'b0000001000;
assign label_1[906] = 10'b0000000100;
assign label_1[907] = 10'b0000001000;
assign label_1[908] = 10'b0000000100;
assign label_1[909] = 10'b0000000100;
assign label_1[910] = 10'b0000000100;
assign label_1[911] = 10'b0000000100;
assign label_1[912] = 10'b0000010000;
assign label_1[913] = 10'b0100000000;
assign label_1[914] = 10'b0100000000;
assign label_1[915] = 10'b0100000000;
assign label_1[916] = 10'b0001000000;
assign label_1[917] = 10'b0001000000;
assign label_1[918] = 10'b0001000000;
assign label_1[919] = 10'b0001000000;
assign label_1[920] = 10'b0000010000;
assign label_1[921] = 10'b0000010000;
assign label_1[922] = 10'b0000000100;
assign label_1[923] = 10'b0100000000;
assign label_1[924] = 10'b0000001000;
assign label_1[925] = 10'b0000001000;
assign label_1[926] = 10'b0100000000;
assign label_1[927] = 10'b0100000000;
assign label_1[928] = 10'b0000000100;
assign label_1[929] = 10'b0001000000;
assign label_1[930] = 10'b0000010000;
assign label_1[931] = 10'b0000001000;
assign label_1[932] = 10'b0000000100;
assign label_1[933] = 10'b0000001000;
assign label_1[934] = 10'b0000001000;
assign label_1[935] = 10'b0000001000;
assign label_1[936] = 10'b0000000100;
assign label_1[937] = 10'b0001000000;
assign label_1[938] = 10'b0000000100;
assign label_1[939] = 10'b0000000100;
assign label_1[940] = 10'b0000000100;
assign label_1[941] = 10'b0000001000;
assign label_1[942] = 10'b0000000100;
assign label_1[943] = 10'b0001000000;
assign label_1[944] = 10'b0000000100;
assign label_1[945] = 10'b0010000000;
assign label_1[946] = 10'b0100000000;
assign label_1[947] = 10'b0100000000;
assign label_1[948] = 10'b0000000001;
assign label_1[949] = 10'b0000000001;
assign label_1[950] = 10'b0001000000;
assign label_1[951] = 10'b0001000000;
assign label_1[952] = 10'b0000000100;
assign label_1[953] = 10'b0000000100;
assign label_1[954] = 10'b0010000000;
assign label_1[955] = 10'b0010000000;
assign label_1[956] = 10'b0001000000;
assign label_1[957] = 10'b0001000000;
assign label_1[958] = 10'b0001000000;
assign label_1[959] = 10'b0001000000;
assign label_1[960] = 10'b0100000000;
assign label_1[961] = 10'b0000010000;
assign label_1[962] = 10'b0100000000;
assign label_1[963] = 10'b1000000000;
assign label_1[964] = 10'b0000010000;
assign label_1[965] = 10'b0000010000;
assign label_1[966] = 10'b1000000000;
assign label_1[967] = 10'b0000010000;
assign label_1[968] = 10'b0000100000;
assign label_1[969] = 10'b0000000001;
assign label_1[970] = 10'b0100000000;
assign label_1[971] = 10'b0100000000;
assign label_1[972] = 10'b0000010000;
assign label_1[973] = 10'b0000001000;
assign label_1[974] = 10'b0100000000;
assign label_1[975] = 10'b0000001000;
assign label_1[976] = 10'b0001000000;
assign label_1[977] = 10'b0000010000;
assign label_1[978] = 10'b0100000000;
assign label_1[979] = 10'b0001000000;
assign label_1[980] = 10'b0000010000;
assign label_1[981] = 10'b0100000000;
assign label_1[982] = 10'b0100000000;
assign label_1[983] = 10'b0000100000;
assign label_1[984] = 10'b0001000000;
assign label_1[985] = 10'b0001000000;
assign label_1[986] = 10'b0001000000;
assign label_1[987] = 10'b0001000000;
assign label_1[988] = 10'b0001000000;
assign label_1[989] = 10'b0001000000;
assign label_1[990] = 10'b0001000000;
assign label_1[991] = 10'b0001000000;
assign label_1[992] = 10'b0001000000;
assign label_1[993] = 10'b0000010000;
assign label_1[994] = 10'b0100000000;
assign label_1[995] = 10'b1000000000;
assign label_1[996] = 10'b0001000000;
assign label_1[997] = 10'b0000000100;
assign label_1[998] = 10'b0001000000;
assign label_1[999] = 10'b0001000000;
assign label_1[1000] = 10'b0000010000;
assign label_1[1001] = 10'b0100000000;
assign label_1[1002] = 10'b0100000000;
assign label_1[1003] = 10'b0001000000;
assign label_1[1004] = 10'b0001000000;
assign label_1[1005] = 10'b0100000000;
assign label_1[1006] = 10'b1000000000;
assign label_1[1007] = 10'b1000000000;
assign label_1[1008] = 10'b0000010000;
assign label_1[1009] = 10'b0000010000;
assign label_1[1010] = 10'b0000000001;
assign label_1[1011] = 10'b0000000001;
assign label_1[1012] = 10'b0000001000;
assign label_1[1013] = 10'b0000001000;
assign label_1[1014] = 10'b0001000000;
assign label_1[1015] = 10'b0001000000;
assign label_1[1016] = 10'b0100000000;
assign label_1[1017] = 10'b0000000100;
assign label_1[1018] = 10'b0100000000;
assign label_1[1019] = 10'b0100000000;
assign label_1[1020] = 10'b0100000000;
assign label_1[1021] = 10'b0000100000;
assign label_1[1022] = 10'b0100000000;
assign label_1[1023] = 10'b0100000000;
assign label_2[0] = 10'b0000100000;
assign label_2[1] = 10'b0000000001;
assign label_2[2] = 10'b0010000000;
assign label_2[3] = 10'b0000100000;
assign label_2[4] = 10'b0010000000;
assign label_2[5] = 10'b0000000100;
assign label_2[6] = 10'b0000000100;
assign label_2[7] = 10'b0000010000;
assign label_2[8] = 10'b0010000000;
assign label_2[9] = 10'b0001000000;
assign label_2[10] = 10'b0000100000;
assign label_2[11] = 10'b0001000000;
assign label_2[12] = 10'b0000001000;
assign label_2[13] = 10'b0001000000;
assign label_2[14] = 10'b1000000000;
assign label_2[15] = 10'b0000010000;
assign label_2[16] = 10'b0000000001;
assign label_2[17] = 10'b0001000000;
assign label_2[18] = 10'b0000000001;
assign label_2[19] = 10'b0000000100;
assign label_2[20] = 10'b0000100000;
assign label_2[21] = 10'b0000000001;
assign label_2[22] = 10'b0000100000;
assign label_2[23] = 10'b0001000000;
assign label_2[24] = 10'b0000000001;
assign label_2[25] = 10'b0000100000;
assign label_2[26] = 10'b0000000001;
assign label_2[27] = 10'b0001000000;
assign label_2[28] = 10'b0001000000;
assign label_2[29] = 10'b0001000000;
assign label_2[30] = 10'b0001000000;
assign label_2[31] = 10'b0001000000;
assign label_2[32] = 10'b0000000010;
assign label_2[33] = 10'b0000100000;
assign label_2[34] = 10'b0000000010;
assign label_2[35] = 10'b0000100000;
assign label_2[36] = 10'b0000000100;
assign label_2[37] = 10'b0001000000;
assign label_2[38] = 10'b0001000000;
assign label_2[39] = 10'b1000000000;
assign label_2[40] = 10'b1000000000;
assign label_2[41] = 10'b0010000000;
assign label_2[42] = 10'b0100000000;
assign label_2[43] = 10'b0000000010;
assign label_2[44] = 10'b0000000100;
assign label_2[45] = 10'b0001000000;
assign label_2[46] = 10'b0001000000;
assign label_2[47] = 10'b0000000001;
assign label_2[48] = 10'b0000001000;
assign label_2[49] = 10'b0000100000;
assign label_2[50] = 10'b0010000000;
assign label_2[51] = 10'b0000000100;
assign label_2[52] = 10'b0000000100;
assign label_2[53] = 10'b0010000000;
assign label_2[54] = 10'b0000010000;
assign label_2[55] = 10'b0000000010;
assign label_2[56] = 10'b1000000000;
assign label_2[57] = 10'b0000001000;
assign label_2[58] = 10'b0000100000;
assign label_2[59] = 10'b0000001000;
assign label_2[60] = 10'b0000000010;
assign label_2[61] = 10'b1000000000;
assign label_2[62] = 10'b0100000000;
assign label_2[63] = 10'b0010000000;
assign label_2[64] = 10'b0010000000;
assign label_2[65] = 10'b0000000100;
assign label_2[66] = 10'b1000000000;
assign label_2[67] = 10'b0000000001;
assign label_2[68] = 10'b0001000000;
assign label_2[69] = 10'b1000000000;
assign label_2[70] = 10'b0010000000;
assign label_2[71] = 10'b0000000001;
assign label_2[72] = 10'b0000001000;
assign label_2[73] = 10'b0001000000;
assign label_2[74] = 10'b0000000100;
assign label_2[75] = 10'b0000010000;
assign label_2[76] = 10'b0000000100;
assign label_2[77] = 10'b0000000100;
assign label_2[78] = 10'b0000000100;
assign label_2[79] = 10'b0000000100;
assign label_2[80] = 10'b0000100000;
assign label_2[81] = 10'b0000000001;
assign label_2[82] = 10'b0000010000;
assign label_2[83] = 10'b0000000100;
assign label_2[84] = 10'b0000100000;
assign label_2[85] = 10'b0000001000;
assign label_2[86] = 10'b0000000001;
assign label_2[87] = 10'b0010000000;
assign label_2[88] = 10'b0010000000;
assign label_2[89] = 10'b0000100000;
assign label_2[90] = 10'b0000000001;
assign label_2[91] = 10'b0000000100;
assign label_2[92] = 10'b0000000100;
assign label_2[93] = 10'b0000000001;
assign label_2[94] = 10'b0000000100;
assign label_2[95] = 10'b0000000001;
assign label_2[96] = 10'b0000000010;
assign label_2[97] = 10'b0000000010;
assign label_2[98] = 10'b1000000000;
assign label_2[99] = 10'b0000001000;
assign label_2[100] = 10'b0000100000;
assign label_2[101] = 10'b0100000000;
assign label_2[102] = 10'b0000001000;
assign label_2[103] = 10'b0100000000;
assign label_2[104] = 10'b0000001000;
assign label_2[105] = 10'b0100000000;
assign label_2[106] = 10'b0000000100;
assign label_2[107] = 10'b0000000100;
assign label_2[108] = 10'b0000000010;
assign label_2[109] = 10'b0100000000;
assign label_2[110] = 10'b0000000010;
assign label_2[111] = 10'b0000000100;
assign label_2[112] = 10'b0000100000;
assign label_2[113] = 10'b0001000000;
assign label_2[114] = 10'b0000001000;
assign label_2[115] = 10'b0000100000;
assign label_2[116] = 10'b0000000100;
assign label_2[117] = 10'b0100000000;
assign label_2[118] = 10'b0100000000;
assign label_2[119] = 10'b0000010000;
assign label_2[120] = 10'b0000001000;
assign label_2[121] = 10'b0100000000;
assign label_2[122] = 10'b0000001000;
assign label_2[123] = 10'b0000100000;
assign label_2[124] = 10'b0010000000;
assign label_2[125] = 10'b0100000000;
assign label_2[126] = 10'b0100000000;
assign label_2[127] = 10'b0000001000;
assign label_2[128] = 10'b0010000000;
assign label_2[129] = 10'b1000000000;
assign label_2[130] = 10'b1000000000;
assign label_2[131] = 10'b0010000000;
assign label_2[132] = 10'b0000000100;
assign label_2[133] = 10'b0000000100;
assign label_2[134] = 10'b0100000000;
assign label_2[135] = 10'b0000001000;
assign label_2[136] = 10'b0000001000;
assign label_2[137] = 10'b0000000100;
assign label_2[138] = 10'b1000000000;
assign label_2[139] = 10'b0010000000;
assign label_2[140] = 10'b1000000000;
assign label_2[141] = 10'b0001000000;
assign label_2[142] = 10'b0000010000;
assign label_2[143] = 10'b0001000000;
assign label_2[144] = 10'b0000100000;
assign label_2[145] = 10'b0000001000;
assign label_2[146] = 10'b0000001000;
assign label_2[147] = 10'b1000000000;
assign label_2[148] = 10'b0000001000;
assign label_2[149] = 10'b0000000100;
assign label_2[150] = 10'b0000100000;
assign label_2[151] = 10'b0000001000;
assign label_2[152] = 10'b0000000100;
assign label_2[153] = 10'b0000000100;
assign label_2[154] = 10'b0000000100;
assign label_2[155] = 10'b0001000000;
assign label_2[156] = 10'b0100000000;
assign label_2[157] = 10'b0100000000;
assign label_2[158] = 10'b0010000000;
assign label_2[159] = 10'b0010000000;
assign label_2[160] = 10'b0010000000;
assign label_2[161] = 10'b0010000000;
assign label_2[162] = 10'b0001000000;
assign label_2[163] = 10'b1000000000;
assign label_2[164] = 10'b1000000000;
assign label_2[165] = 10'b0000010000;
assign label_2[166] = 10'b0000010000;
assign label_2[167] = 10'b1000000000;
assign label_2[168] = 10'b0010000000;
assign label_2[169] = 10'b1000000000;
assign label_2[170] = 10'b0010000000;
assign label_2[171] = 10'b0000001000;
assign label_2[172] = 10'b0000010000;
assign label_2[173] = 10'b0000010000;
assign label_2[174] = 10'b0000001000;
assign label_2[175] = 10'b1000000000;
assign label_2[176] = 10'b1000000000;
assign label_2[177] = 10'b0001000000;
assign label_2[178] = 10'b0000010000;
assign label_2[179] = 10'b0000100000;
assign label_2[180] = 10'b0001000000;
assign label_2[181] = 10'b0001000000;
assign label_2[182] = 10'b0000001000;
assign label_2[183] = 10'b0001000000;
assign label_2[184] = 10'b0000010000;
assign label_2[185] = 10'b0000001000;
assign label_2[186] = 10'b0010000000;
assign label_2[187] = 10'b0000000001;
assign label_2[188] = 10'b0010000000;
assign label_2[189] = 10'b0000010000;
assign label_2[190] = 10'b0000010000;
assign label_2[191] = 10'b1000000000;
assign label_2[192] = 10'b0000010000;
assign label_2[193] = 10'b0000001000;
assign label_2[194] = 10'b0000010000;
assign label_2[195] = 10'b0000100000;
assign label_2[196] = 10'b0000100000;
assign label_2[197] = 10'b0100000000;
assign label_2[198] = 10'b0000001000;
assign label_2[199] = 10'b1000000000;
assign label_2[200] = 10'b0000010000;
assign label_2[201] = 10'b0010000000;
assign label_2[202] = 10'b0000000100;
assign label_2[203] = 10'b0100000000;
assign label_2[204] = 10'b0000000100;
assign label_2[205] = 10'b0000001000;
assign label_2[206] = 10'b0100000000;
assign label_2[207] = 10'b0100000000;
assign label_2[208] = 10'b0000000100;
assign label_2[209] = 10'b0000010000;
assign label_2[210] = 10'b0000010000;
assign label_2[211] = 10'b0100000000;
assign label_2[212] = 10'b0100000000;
assign label_2[213] = 10'b0100000000;
assign label_2[214] = 10'b0000001000;
assign label_2[215] = 10'b0100000000;
assign label_2[216] = 10'b0000000100;
assign label_2[217] = 10'b0000000100;
assign label_2[218] = 10'b0000010000;
assign label_2[219] = 10'b0000100000;
assign label_2[220] = 10'b0001000000;
assign label_2[221] = 10'b0001000000;
assign label_2[222] = 10'b0001000000;
assign label_2[223] = 10'b0001000000;
assign label_2[224] = 10'b0000001000;
assign label_2[225] = 10'b1000000000;
assign label_2[226] = 10'b0000100000;
assign label_2[227] = 10'b0000001000;
assign label_2[228] = 10'b0001000000;
assign label_2[229] = 10'b0001000000;
assign label_2[230] = 10'b1000000000;
assign label_2[231] = 10'b0001000000;
assign label_2[232] = 10'b0000001000;
assign label_2[233] = 10'b0000100000;
assign label_2[234] = 10'b0010000000;
assign label_2[235] = 10'b1000000000;
assign label_2[236] = 10'b0000001000;
assign label_2[237] = 10'b0100000000;
assign label_2[238] = 10'b0000001000;
assign label_2[239] = 10'b0100000000;
assign label_2[240] = 10'b1000000000;
assign label_2[241] = 10'b1000000000;
assign label_2[242] = 10'b0000000100;
assign label_2[243] = 10'b0000000100;
assign label_2[244] = 10'b0000100000;
assign label_2[245] = 10'b0100000000;
assign label_2[246] = 10'b0000001000;
assign label_2[247] = 10'b1000000000;
assign label_2[248] = 10'b1000000000;
assign label_2[249] = 10'b0100000000;
assign label_2[250] = 10'b0010000000;
assign label_2[251] = 10'b0001000000;
assign label_2[252] = 10'b0000000100;
assign label_2[253] = 10'b0100000000;
assign label_2[254] = 10'b0000000100;
assign label_2[255] = 10'b0001000000;
assign label_2[256] = 10'b0000010000;
assign label_2[257] = 10'b0001000000;
assign label_2[258] = 10'b0000001000;
assign label_2[259] = 10'b0000010000;
assign label_2[260] = 10'b0000010000;
assign label_2[261] = 10'b0000100000;
assign label_2[262] = 10'b0000001000;
assign label_2[263] = 10'b0001000000;
assign label_2[264] = 10'b0000010000;
assign label_2[265] = 10'b0000010000;
assign label_2[266] = 10'b0000010000;
assign label_2[267] = 10'b0000010000;
assign label_2[268] = 10'b0000010000;
assign label_2[269] = 10'b0010000000;
assign label_2[270] = 10'b0001000000;
assign label_2[271] = 10'b0001000000;
assign label_2[272] = 10'b0000001000;
assign label_2[273] = 10'b0000100000;
assign label_2[274] = 10'b0000000100;
assign label_2[275] = 10'b0000000100;
assign label_2[276] = 10'b0000000100;
assign label_2[277] = 10'b0000000100;
assign label_2[278] = 10'b0000000100;
assign label_2[279] = 10'b0000000100;
assign label_2[280] = 10'b0000010000;
assign label_2[281] = 10'b0000000001;
assign label_2[282] = 10'b0000100000;
assign label_2[283] = 10'b0000000100;
assign label_2[284] = 10'b0001000000;
assign label_2[285] = 10'b0000000001;
assign label_2[286] = 10'b0000100000;
assign label_2[287] = 10'b0001000000;
assign label_2[288] = 10'b0001000000;
assign label_2[289] = 10'b0000010000;
assign label_2[290] = 10'b0001000000;
assign label_2[291] = 10'b0000010000;
assign label_2[292] = 10'b0100000000;
assign label_2[293] = 10'b0000100000;
assign label_2[294] = 10'b0000100000;
assign label_2[295] = 10'b0000000001;
assign label_2[296] = 10'b0001000000;
assign label_2[297] = 10'b0000010000;
assign label_2[298] = 10'b0000000100;
assign label_2[299] = 10'b0000010000;
assign label_2[300] = 10'b0000010000;
assign label_2[301] = 10'b1000000000;
assign label_2[302] = 10'b0000010000;
assign label_2[303] = 10'b0000010000;
assign label_2[304] = 10'b0000010000;
assign label_2[305] = 10'b0000010000;
assign label_2[306] = 10'b0000000001;
assign label_2[307] = 10'b0000010000;
assign label_2[308] = 10'b0000000100;
assign label_2[309] = 10'b0000010000;
assign label_2[310] = 10'b0000000010;
assign label_2[311] = 10'b0000100000;
assign label_2[312] = 10'b0000100000;
assign label_2[313] = 10'b0000000001;
assign label_2[314] = 10'b0000010000;
assign label_2[315] = 10'b0001000000;
assign label_2[316] = 10'b0001000000;
assign label_2[317] = 10'b0001000000;
assign label_2[318] = 10'b0000000100;
assign label_2[319] = 10'b0000010000;
assign label_2[320] = 10'b0000000100;
assign label_2[321] = 10'b0000000100;
assign label_2[322] = 10'b0001000000;
assign label_2[323] = 10'b0001000000;
assign label_2[324] = 10'b0000100000;
assign label_2[325] = 10'b0000010000;
assign label_2[326] = 10'b0000010000;
assign label_2[327] = 10'b0001000000;
assign label_2[328] = 10'b0000001000;
assign label_2[329] = 10'b0000001000;
assign label_2[330] = 10'b0000100000;
assign label_2[331] = 10'b0100000000;
assign label_2[332] = 10'b0100000000;
assign label_2[333] = 10'b0000000001;
assign label_2[334] = 10'b0000100000;
assign label_2[335] = 10'b0100000000;
assign label_2[336] = 10'b0000000100;
assign label_2[337] = 10'b0000000100;
assign label_2[338] = 10'b0100000000;
assign label_2[339] = 10'b0100000000;
assign label_2[340] = 10'b0000000100;
assign label_2[341] = 10'b0000000100;
assign label_2[342] = 10'b0000000100;
assign label_2[343] = 10'b0000000100;
assign label_2[344] = 10'b0000001000;
assign label_2[345] = 10'b0000001000;
assign label_2[346] = 10'b0000000100;
assign label_2[347] = 10'b0000000100;
assign label_2[348] = 10'b0000000100;
assign label_2[349] = 10'b0000000100;
assign label_2[350] = 10'b0000000100;
assign label_2[351] = 10'b0000000100;
assign label_2[352] = 10'b0000010000;
assign label_2[353] = 10'b0001000000;
assign label_2[354] = 10'b0000010000;
assign label_2[355] = 10'b0000000100;
assign label_2[356] = 10'b0000000100;
assign label_2[357] = 10'b0000010000;
assign label_2[358] = 10'b1000000000;
assign label_2[359] = 10'b0001000000;
assign label_2[360] = 10'b0100000000;
assign label_2[361] = 10'b0000100000;
assign label_2[362] = 10'b0000000001;
assign label_2[363] = 10'b0000010000;
assign label_2[364] = 10'b0000100000;
assign label_2[365] = 10'b0000100000;
assign label_2[366] = 10'b0001000000;
assign label_2[367] = 10'b0001000000;
assign label_2[368] = 10'b0000000001;
assign label_2[369] = 10'b0000000001;
assign label_2[370] = 10'b0100000000;
assign label_2[371] = 10'b0001000000;
assign label_2[372] = 10'b0000100000;
assign label_2[373] = 10'b0001000000;
assign label_2[374] = 10'b0001000000;
assign label_2[375] = 10'b0000000100;
assign label_2[376] = 10'b0000100000;
assign label_2[377] = 10'b0000100000;
assign label_2[378] = 10'b0100000000;
assign label_2[379] = 10'b0100000000;
assign label_2[380] = 10'b0000001000;
assign label_2[381] = 10'b0100000000;
assign label_2[382] = 10'b0001000000;
assign label_2[383] = 10'b0100000000;
assign label_2[384] = 10'b1000000000;
assign label_2[385] = 10'b0000010000;
assign label_2[386] = 10'b1000000000;
assign label_2[387] = 10'b0000010000;
assign label_2[388] = 10'b1000000000;
assign label_2[389] = 10'b0000100000;
assign label_2[390] = 10'b1000000000;
assign label_2[391] = 10'b0000000100;
assign label_2[392] = 10'b1000000000;
assign label_2[393] = 10'b1000000000;
assign label_2[394] = 10'b0010000000;
assign label_2[395] = 10'b0000000100;
assign label_2[396] = 10'b0000100000;
assign label_2[397] = 10'b0000100000;
assign label_2[398] = 10'b1000000000;
assign label_2[399] = 10'b0000000100;
assign label_2[400] = 10'b0000100000;
assign label_2[401] = 10'b0000000100;
assign label_2[402] = 10'b0000010000;
assign label_2[403] = 10'b0000100000;
assign label_2[404] = 10'b0000001000;
assign label_2[405] = 10'b0000010000;
assign label_2[406] = 10'b1000000000;
assign label_2[407] = 10'b0000001000;
assign label_2[408] = 10'b0000010000;
assign label_2[409] = 10'b0000001000;
assign label_2[410] = 10'b1000000000;
assign label_2[411] = 10'b0000100000;
assign label_2[412] = 10'b0000001000;
assign label_2[413] = 10'b0000001000;
assign label_2[414] = 10'b0000001000;
assign label_2[415] = 10'b0100000000;
assign label_2[416] = 10'b0000010000;
assign label_2[417] = 10'b1000000000;
assign label_2[418] = 10'b0001000000;
assign label_2[419] = 10'b0000000100;
assign label_2[420] = 10'b0001000000;
assign label_2[421] = 10'b0000000100;
assign label_2[422] = 10'b0000000001;
assign label_2[423] = 10'b0000000100;
assign label_2[424] = 10'b0001000000;
assign label_2[425] = 10'b0000000100;
assign label_2[426] = 10'b0001000000;
assign label_2[427] = 10'b0000000100;
assign label_2[428] = 10'b0000010000;
assign label_2[429] = 10'b0000000100;
assign label_2[430] = 10'b0000000100;
assign label_2[431] = 10'b0000000100;
assign label_2[432] = 10'b0000000001;
assign label_2[433] = 10'b0001000000;
assign label_2[434] = 10'b0000100000;
assign label_2[435] = 10'b0000001000;
assign label_2[436] = 10'b0100000000;
assign label_2[437] = 10'b0100000000;
assign label_2[438] = 10'b0100000000;
assign label_2[439] = 10'b0000001000;
assign label_2[440] = 10'b0000000001;
assign label_2[441] = 10'b1000000000;
assign label_2[442] = 10'b0100000000;
assign label_2[443] = 10'b0001000000;
assign label_2[444] = 10'b0001000000;
assign label_2[445] = 10'b0000000001;
assign label_2[446] = 10'b0100000000;
assign label_2[447] = 10'b0100000000;
assign label_2[448] = 10'b0001000000;
assign label_2[449] = 10'b0000010000;
assign label_2[450] = 10'b0000100000;
assign label_2[451] = 10'b0000100000;
assign label_2[452] = 10'b0001000000;
assign label_2[453] = 10'b0001000000;
assign label_2[454] = 10'b0000000001;
assign label_2[455] = 10'b0000000001;
assign label_2[456] = 10'b0001000000;
assign label_2[457] = 10'b0001000000;
assign label_2[458] = 10'b0001000000;
assign label_2[459] = 10'b0000000100;
assign label_2[460] = 10'b0001000000;
assign label_2[461] = 10'b0001000000;
assign label_2[462] = 10'b0100000000;
assign label_2[463] = 10'b0100000000;
assign label_2[464] = 10'b0001000000;
assign label_2[465] = 10'b0001000000;
assign label_2[466] = 10'b0000000100;
assign label_2[467] = 10'b0000000100;
assign label_2[468] = 10'b0000000100;
assign label_2[469] = 10'b0000000100;
assign label_2[470] = 10'b0000000100;
assign label_2[471] = 10'b0000000100;
assign label_2[472] = 10'b0001000000;
assign label_2[473] = 10'b0001000000;
assign label_2[474] = 10'b0001000000;
assign label_2[475] = 10'b0001000000;
assign label_2[476] = 10'b0000000001;
assign label_2[477] = 10'b0000000001;
assign label_2[478] = 10'b0000000100;
assign label_2[479] = 10'b0000000100;
assign label_2[480] = 10'b0000000100;
assign label_2[481] = 10'b0000000100;
assign label_2[482] = 10'b0000000100;
assign label_2[483] = 10'b0000000100;
assign label_2[484] = 10'b0000000100;
assign label_2[485] = 10'b0000000100;
assign label_2[486] = 10'b0000000100;
assign label_2[487] = 10'b0000000100;
assign label_2[488] = 10'b0000000100;
assign label_2[489] = 10'b0000000100;
assign label_2[490] = 10'b0000000100;
assign label_2[491] = 10'b0000000100;
assign label_2[492] = 10'b0000000100;
assign label_2[493] = 10'b0000000100;
assign label_2[494] = 10'b0000000100;
assign label_2[495] = 10'b0000000100;
assign label_2[496] = 10'b0000000100;
assign label_2[497] = 10'b0000000100;
assign label_2[498] = 10'b0000000100;
assign label_2[499] = 10'b0000000100;
assign label_2[500] = 10'b0000000100;
assign label_2[501] = 10'b0000000100;
assign label_2[502] = 10'b0000000100;
assign label_2[503] = 10'b0000000100;
assign label_2[504] = 10'b0000000100;
assign label_2[505] = 10'b0000000100;
assign label_2[506] = 10'b0000000100;
assign label_2[507] = 10'b0000000100;
assign label_2[508] = 10'b0000000100;
assign label_2[509] = 10'b0000000100;
assign label_2[510] = 10'b0000000100;
assign label_2[511] = 10'b0000000100;
assign label_2[512] = 10'b0000001000;
assign label_2[513] = 10'b0000001000;
assign label_2[514] = 10'b0000001000;
assign label_2[515] = 10'b0000100000;
assign label_2[516] = 10'b0000001000;
assign label_2[517] = 10'b0000100000;
assign label_2[518] = 10'b0000000100;
assign label_2[519] = 10'b0000000100;
assign label_2[520] = 10'b0000000010;
assign label_2[521] = 10'b0000100000;
assign label_2[522] = 10'b0000000100;
assign label_2[523] = 10'b0000000001;
assign label_2[524] = 10'b0000000010;
assign label_2[525] = 10'b0000100000;
assign label_2[526] = 10'b0000000100;
assign label_2[527] = 10'b0000100000;
assign label_2[528] = 10'b0000100000;
assign label_2[529] = 10'b0000000100;
assign label_2[530] = 10'b0000000100;
assign label_2[531] = 10'b0000000100;
assign label_2[532] = 10'b0000001000;
assign label_2[533] = 10'b0000000100;
assign label_2[534] = 10'b0000000100;
assign label_2[535] = 10'b0000000100;
assign label_2[536] = 10'b0001000000;
assign label_2[537] = 10'b0000000001;
assign label_2[538] = 10'b0000000001;
assign label_2[539] = 10'b0000100000;
assign label_2[540] = 10'b0000000001;
assign label_2[541] = 10'b0000000100;
assign label_2[542] = 10'b0000000100;
assign label_2[543] = 10'b0000000001;
assign label_2[544] = 10'b0000000001;
assign label_2[545] = 10'b0000100000;
assign label_2[546] = 10'b0000000001;
assign label_2[547] = 10'b0000001000;
assign label_2[548] = 10'b0000000001;
assign label_2[549] = 10'b0000100000;
assign label_2[550] = 10'b0000100000;
assign label_2[551] = 10'b0000100000;
assign label_2[552] = 10'b0000000001;
assign label_2[553] = 10'b0000000001;
assign label_2[554] = 10'b0000000001;
assign label_2[555] = 10'b0000000001;
assign label_2[556] = 10'b0000100000;
assign label_2[557] = 10'b0000100000;
assign label_2[558] = 10'b0000100000;
assign label_2[559] = 10'b0000100000;
assign label_2[560] = 10'b0000100000;
assign label_2[561] = 10'b0000100000;
assign label_2[562] = 10'b0000001000;
assign label_2[563] = 10'b0000001000;
assign label_2[564] = 10'b0000000100;
assign label_2[565] = 10'b0100000000;
assign label_2[566] = 10'b0000100000;
assign label_2[567] = 10'b0000000001;
assign label_2[568] = 10'b0000001000;
assign label_2[569] = 10'b0000001000;
assign label_2[570] = 10'b0000001000;
assign label_2[571] = 10'b0000001000;
assign label_2[572] = 10'b0000000100;
assign label_2[573] = 10'b0000000100;
assign label_2[574] = 10'b0000000100;
assign label_2[575] = 10'b0000000100;
assign label_2[576] = 10'b0000000001;
assign label_2[577] = 10'b0000000001;
assign label_2[578] = 10'b0000000100;
assign label_2[579] = 10'b0000000001;
assign label_2[580] = 10'b0000100000;
assign label_2[581] = 10'b0000100000;
assign label_2[582] = 10'b0000001000;
assign label_2[583] = 10'b0000000100;
assign label_2[584] = 10'b0000000001;
assign label_2[585] = 10'b0000000001;
assign label_2[586] = 10'b0000000001;
assign label_2[587] = 10'b0000000001;
assign label_2[588] = 10'b0000000001;
assign label_2[589] = 10'b0000000100;
assign label_2[590] = 10'b0000000001;
assign label_2[591] = 10'b0000000001;
assign label_2[592] = 10'b0000100000;
assign label_2[593] = 10'b0100000000;
assign label_2[594] = 10'b0000000001;
assign label_2[595] = 10'b0000000001;
assign label_2[596] = 10'b0100000000;
assign label_2[597] = 10'b0100000000;
assign label_2[598] = 10'b0100000000;
assign label_2[599] = 10'b0100000000;
assign label_2[600] = 10'b1000000000;
assign label_2[601] = 10'b1000000000;
assign label_2[602] = 10'b0000000001;
assign label_2[603] = 10'b0000000100;
assign label_2[604] = 10'b0000000010;
assign label_2[605] = 10'b0000000001;
assign label_2[606] = 10'b0100000000;
assign label_2[607] = 10'b0100000000;
assign label_2[608] = 10'b0000000001;
assign label_2[609] = 10'b0000001000;
assign label_2[610] = 10'b0000000100;
assign label_2[611] = 10'b0000000100;
assign label_2[612] = 10'b0000000100;
assign label_2[613] = 10'b0000100000;
assign label_2[614] = 10'b0000000001;
assign label_2[615] = 10'b0000000001;
assign label_2[616] = 10'b0000000001;
assign label_2[617] = 10'b0000000001;
assign label_2[618] = 10'b0000000001;
assign label_2[619] = 10'b0000000001;
assign label_2[620] = 10'b0000000001;
assign label_2[621] = 10'b0000000001;
assign label_2[622] = 10'b0000100000;
assign label_2[623] = 10'b0000000001;
assign label_2[624] = 10'b0000000001;
assign label_2[625] = 10'b0000000001;
assign label_2[626] = 10'b0000000100;
assign label_2[627] = 10'b0001000000;
assign label_2[628] = 10'b0000100000;
assign label_2[629] = 10'b0000100000;
assign label_2[630] = 10'b0100000000;
assign label_2[631] = 10'b0000100000;
assign label_2[632] = 10'b0000100000;
assign label_2[633] = 10'b0000100000;
assign label_2[634] = 10'b0000000100;
assign label_2[635] = 10'b0000000001;
assign label_2[636] = 10'b0000000100;
assign label_2[637] = 10'b0000000001;
assign label_2[638] = 10'b0000000001;
assign label_2[639] = 10'b0000000001;
assign label_2[640] = 10'b0000100000;
assign label_2[641] = 10'b0000000001;
assign label_2[642] = 10'b0000100000;
assign label_2[643] = 10'b0100000000;
assign label_2[644] = 10'b0000100000;
assign label_2[645] = 10'b0000100000;
assign label_2[646] = 10'b0001000000;
assign label_2[647] = 10'b0001000000;
assign label_2[648] = 10'b0000001000;
assign label_2[649] = 10'b0000000100;
assign label_2[650] = 10'b0000000100;
assign label_2[651] = 10'b0100000000;
assign label_2[652] = 10'b0000000001;
assign label_2[653] = 10'b0000100000;
assign label_2[654] = 10'b0000000100;
assign label_2[655] = 10'b0000000100;
assign label_2[656] = 10'b0000001000;
assign label_2[657] = 10'b0100000000;
assign label_2[658] = 10'b0000001000;
assign label_2[659] = 10'b0000000010;
assign label_2[660] = 10'b0000000100;
assign label_2[661] = 10'b0100000000;
assign label_2[662] = 10'b0000000010;
assign label_2[663] = 10'b0001000000;
assign label_2[664] = 10'b0100000000;
assign label_2[665] = 10'b0000100000;
assign label_2[666] = 10'b0000100000;
assign label_2[667] = 10'b0000100000;
assign label_2[668] = 10'b0000100000;
assign label_2[669] = 10'b0100000000;
assign label_2[670] = 10'b0000000100;
assign label_2[671] = 10'b0000001000;
assign label_2[672] = 10'b0000000100;
assign label_2[673] = 10'b1000000000;
assign label_2[674] = 10'b0010000000;
assign label_2[675] = 10'b0100000000;
assign label_2[676] = 10'b0000000100;
assign label_2[677] = 10'b0000000100;
assign label_2[678] = 10'b0000000100;
assign label_2[679] = 10'b0100000000;
assign label_2[680] = 10'b0010000000;
assign label_2[681] = 10'b0000000100;
assign label_2[682] = 10'b0000000100;
assign label_2[683] = 10'b0000000100;
assign label_2[684] = 10'b0100000000;
assign label_2[685] = 10'b0000000100;
assign label_2[686] = 10'b0100000000;
assign label_2[687] = 10'b0100000000;
assign label_2[688] = 10'b0000000001;
assign label_2[689] = 10'b0010000000;
assign label_2[690] = 10'b0000000100;
assign label_2[691] = 10'b0000000001;
assign label_2[692] = 10'b0100000000;
assign label_2[693] = 10'b0000010000;
assign label_2[694] = 10'b0000000100;
assign label_2[695] = 10'b0100000000;
assign label_2[696] = 10'b0100000000;
assign label_2[697] = 10'b0000000001;
assign label_2[698] = 10'b0000000100;
assign label_2[699] = 10'b0000000100;
assign label_2[700] = 10'b0000000001;
assign label_2[701] = 10'b0100000000;
assign label_2[702] = 10'b0000000100;
assign label_2[703] = 10'b0000000100;
assign label_2[704] = 10'b0010000000;
assign label_2[705] = 10'b0000000100;
assign label_2[706] = 10'b0001000000;
assign label_2[707] = 10'b0000000001;
assign label_2[708] = 10'b0010000000;
assign label_2[709] = 10'b0010000000;
assign label_2[710] = 10'b0010000000;
assign label_2[711] = 10'b0100000000;
assign label_2[712] = 10'b0000000100;
assign label_2[713] = 10'b0001000000;
assign label_2[714] = 10'b0000000100;
assign label_2[715] = 10'b0000000100;
assign label_2[716] = 10'b0000001000;
assign label_2[717] = 10'b0000001000;
assign label_2[718] = 10'b0100000000;
assign label_2[719] = 10'b0100000000;
assign label_2[720] = 10'b0000000100;
assign label_2[721] = 10'b0000000100;
assign label_2[722] = 10'b0000000100;
assign label_2[723] = 10'b0100000000;
assign label_2[724] = 10'b0010000000;
assign label_2[725] = 10'b0010000000;
assign label_2[726] = 10'b0000000100;
assign label_2[727] = 10'b0000000100;
assign label_2[728] = 10'b0000001000;
assign label_2[729] = 10'b0000001000;
assign label_2[730] = 10'b0000001000;
assign label_2[731] = 10'b0000001000;
assign label_2[732] = 10'b0100000000;
assign label_2[733] = 10'b0100000000;
assign label_2[734] = 10'b0100000000;
assign label_2[735] = 10'b0100000000;
assign label_2[736] = 10'b0010000000;
assign label_2[737] = 10'b0000000001;
assign label_2[738] = 10'b0001000000;
assign label_2[739] = 10'b0010000000;
assign label_2[740] = 10'b0010000000;
assign label_2[741] = 10'b0000000001;
assign label_2[742] = 10'b0100000000;
assign label_2[743] = 10'b0000000100;
assign label_2[744] = 10'b0100000000;
assign label_2[745] = 10'b0100000000;
assign label_2[746] = 10'b0000010000;
assign label_2[747] = 10'b1000000000;
assign label_2[748] = 10'b0000000100;
assign label_2[749] = 10'b0000000001;
assign label_2[750] = 10'b0000100000;
assign label_2[751] = 10'b0001000000;
assign label_2[752] = 10'b0000000001;
assign label_2[753] = 10'b0000000001;
assign label_2[754] = 10'b0000000100;
assign label_2[755] = 10'b0000000100;
assign label_2[756] = 10'b0001000000;
assign label_2[757] = 10'b0001000000;
assign label_2[758] = 10'b0000000100;
assign label_2[759] = 10'b0000000100;
assign label_2[760] = 10'b0001000000;
assign label_2[761] = 10'b0100000000;
assign label_2[762] = 10'b0000000001;
assign label_2[763] = 10'b0000000100;
assign label_2[764] = 10'b0000010000;
assign label_2[765] = 10'b0000000100;
assign label_2[766] = 10'b0000000001;
assign label_2[767] = 10'b0000000100;
assign label_2[768] = 10'b0000100000;
assign label_2[769] = 10'b0000100000;
assign label_2[770] = 10'b0000000100;
assign label_2[771] = 10'b0000001000;
assign label_2[772] = 10'b0000001000;
assign label_2[773] = 10'b0000001000;
assign label_2[774] = 10'b0000100000;
assign label_2[775] = 10'b0000001000;
assign label_2[776] = 10'b0000100000;
assign label_2[777] = 10'b0000001000;
assign label_2[778] = 10'b0000001000;
assign label_2[779] = 10'b0000000010;
assign label_2[780] = 10'b0000000100;
assign label_2[781] = 10'b0000100000;
assign label_2[782] = 10'b0000001000;
assign label_2[783] = 10'b0000000100;
assign label_2[784] = 10'b0000100000;
assign label_2[785] = 10'b0000100000;
assign label_2[786] = 10'b0000001000;
assign label_2[787] = 10'b0000001000;
assign label_2[788] = 10'b0000100000;
assign label_2[789] = 10'b0100000000;
assign label_2[790] = 10'b0000100000;
assign label_2[791] = 10'b0000001000;
assign label_2[792] = 10'b0000100000;
assign label_2[793] = 10'b0010000000;
assign label_2[794] = 10'b0100000000;
assign label_2[795] = 10'b0000001000;
assign label_2[796] = 10'b0000100000;
assign label_2[797] = 10'b1000000000;
assign label_2[798] = 10'b0000100000;
assign label_2[799] = 10'b0100000000;
assign label_2[800] = 10'b0000001000;
assign label_2[801] = 10'b0000100000;
assign label_2[802] = 10'b0000100000;
assign label_2[803] = 10'b0001000000;
assign label_2[804] = 10'b0000100000;
assign label_2[805] = 10'b0000000001;
assign label_2[806] = 10'b0001000000;
assign label_2[807] = 10'b0001000000;
assign label_2[808] = 10'b0000001000;
assign label_2[809] = 10'b0000000001;
assign label_2[810] = 10'b0000001000;
assign label_2[811] = 10'b0000100000;
assign label_2[812] = 10'b0100000000;
assign label_2[813] = 10'b0100000000;
assign label_2[814] = 10'b0001000000;
assign label_2[815] = 10'b0000000100;
assign label_2[816] = 10'b0000000001;
assign label_2[817] = 10'b0000000100;
assign label_2[818] = 10'b0000001000;
assign label_2[819] = 10'b0000001000;
assign label_2[820] = 10'b0000100000;
assign label_2[821] = 10'b0000100000;
assign label_2[822] = 10'b0000100000;
assign label_2[823] = 10'b0000100000;
assign label_2[824] = 10'b0000000001;
assign label_2[825] = 10'b0000000100;
assign label_2[826] = 10'b0100000000;
assign label_2[827] = 10'b0000001000;
assign label_2[828] = 10'b0000000100;
assign label_2[829] = 10'b0100000000;
assign label_2[830] = 10'b0001000000;
assign label_2[831] = 10'b0000000100;
assign label_2[832] = 10'b0010000000;
assign label_2[833] = 10'b0000000010;
assign label_2[834] = 10'b0000000100;
assign label_2[835] = 10'b0000000100;
assign label_2[836] = 10'b0000000100;
assign label_2[837] = 10'b0000001000;
assign label_2[838] = 10'b0001000000;
assign label_2[839] = 10'b0001000000;
assign label_2[840] = 10'b0000010000;
assign label_2[841] = 10'b0000000100;
assign label_2[842] = 10'b0000010000;
assign label_2[843] = 10'b1000000000;
assign label_2[844] = 10'b0000001000;
assign label_2[845] = 10'b0000000100;
assign label_2[846] = 10'b0000010000;
assign label_2[847] = 10'b0000000100;
assign label_2[848] = 10'b0000000100;
assign label_2[849] = 10'b0000001000;
assign label_2[850] = 10'b0001000000;
assign label_2[851] = 10'b0000001000;
assign label_2[852] = 10'b0001000000;
assign label_2[853] = 10'b0001000000;
assign label_2[854] = 10'b0000000001;
assign label_2[855] = 10'b0000000100;
assign label_2[856] = 10'b0000000100;
assign label_2[857] = 10'b0000000100;
assign label_2[858] = 10'b0000000100;
assign label_2[859] = 10'b0001000000;
assign label_2[860] = 10'b0100000000;
assign label_2[861] = 10'b0000000100;
assign label_2[862] = 10'b0000000100;
assign label_2[863] = 10'b0000000001;
assign label_2[864] = 10'b0010000000;
assign label_2[865] = 10'b0000010000;
assign label_2[866] = 10'b0010000000;
assign label_2[867] = 10'b0010000000;
assign label_2[868] = 10'b1000000000;
assign label_2[869] = 10'b0010000000;
assign label_2[870] = 10'b1000000000;
assign label_2[871] = 10'b1000000000;
assign label_2[872] = 10'b0010000000;
assign label_2[873] = 10'b0010000000;
assign label_2[874] = 10'b0010000000;
assign label_2[875] = 10'b0010000000;
assign label_2[876] = 10'b1000000000;
assign label_2[877] = 10'b1000000000;
assign label_2[878] = 10'b1000000000;
assign label_2[879] = 10'b1000000000;
assign label_2[880] = 10'b0000010000;
assign label_2[881] = 10'b0000010000;
assign label_2[882] = 10'b0000010000;
assign label_2[883] = 10'b1000000000;
assign label_2[884] = 10'b0010000000;
assign label_2[885] = 10'b0010000000;
assign label_2[886] = 10'b0010000000;
assign label_2[887] = 10'b1000000000;
assign label_2[888] = 10'b0010000000;
assign label_2[889] = 10'b1000000000;
assign label_2[890] = 10'b1000000000;
assign label_2[891] = 10'b1000000000;
assign label_2[892] = 10'b0000010000;
assign label_2[893] = 10'b1000000000;
assign label_2[894] = 10'b0100000000;
assign label_2[895] = 10'b0000010000;
assign label_2[896] = 10'b0000000010;
assign label_2[897] = 10'b0000010000;
assign label_2[898] = 10'b0010000000;
assign label_2[899] = 10'b0100000000;
assign label_2[900] = 10'b1000000000;
assign label_2[901] = 10'b0000010000;
assign label_2[902] = 10'b0010000000;
assign label_2[903] = 10'b0100000000;
assign label_2[904] = 10'b0010000000;
assign label_2[905] = 10'b0000010000;
assign label_2[906] = 10'b0000010000;
assign label_2[907] = 10'b0010000000;
assign label_2[908] = 10'b0010000000;
assign label_2[909] = 10'b0000000100;
assign label_2[910] = 10'b0100000000;
assign label_2[911] = 10'b0000000010;
assign label_2[912] = 10'b0000000100;
assign label_2[913] = 10'b0000000100;
assign label_2[914] = 10'b0000000100;
assign label_2[915] = 10'b0000000100;
assign label_2[916] = 10'b0000000100;
assign label_2[917] = 10'b0000000100;
assign label_2[918] = 10'b0000000100;
assign label_2[919] = 10'b0000000100;
assign label_2[920] = 10'b0100000000;
assign label_2[921] = 10'b1000000000;
assign label_2[922] = 10'b0100000000;
assign label_2[923] = 10'b0100000000;
assign label_2[924] = 10'b0000000100;
assign label_2[925] = 10'b0000000100;
assign label_2[926] = 10'b0000000100;
assign label_2[927] = 10'b0000000100;
assign label_2[928] = 10'b0000000100;
assign label_2[929] = 10'b0100000000;
assign label_2[930] = 10'b0100000000;
assign label_2[931] = 10'b0100000000;
assign label_2[932] = 10'b0001000000;
assign label_2[933] = 10'b0001000000;
assign label_2[934] = 10'b0000000100;
assign label_2[935] = 10'b0100000000;
assign label_2[936] = 10'b0000000100;
assign label_2[937] = 10'b0000000100;
assign label_2[938] = 10'b0001000000;
assign label_2[939] = 10'b0000000100;
assign label_2[940] = 10'b0000001000;
assign label_2[941] = 10'b0000000100;
assign label_2[942] = 10'b0100000000;
assign label_2[943] = 10'b0100000000;
assign label_2[944] = 10'b0000000100;
assign label_2[945] = 10'b0000001000;
assign label_2[946] = 10'b0000001000;
assign label_2[947] = 10'b0000100000;
assign label_2[948] = 10'b0000000100;
assign label_2[949] = 10'b0000000100;
assign label_2[950] = 10'b0000000100;
assign label_2[951] = 10'b0000000100;
assign label_2[952] = 10'b0000000001;
assign label_2[953] = 10'b0000000001;
assign label_2[954] = 10'b0000000001;
assign label_2[955] = 10'b0000000001;
assign label_2[956] = 10'b0000000100;
assign label_2[957] = 10'b0000000001;
assign label_2[958] = 10'b0001000000;
assign label_2[959] = 10'b0100000000;
assign label_2[960] = 10'b0100000000;
assign label_2[961] = 10'b0001000000;
assign label_2[962] = 10'b0000100000;
assign label_2[963] = 10'b0000001000;
assign label_2[964] = 10'b0010000000;
assign label_2[965] = 10'b0010000000;
assign label_2[966] = 10'b0000010000;
assign label_2[967] = 10'b0000000100;
assign label_2[968] = 10'b0100000000;
assign label_2[969] = 10'b0000000100;
assign label_2[970] = 10'b1000000000;
assign label_2[971] = 10'b0000010000;
assign label_2[972] = 10'b0000001000;
assign label_2[973] = 10'b0000100000;
assign label_2[974] = 10'b0100000000;
assign label_2[975] = 10'b0100000000;
assign label_2[976] = 10'b0000010000;
assign label_2[977] = 10'b0100000000;
assign label_2[978] = 10'b0100000000;
assign label_2[979] = 10'b0100000000;
assign label_2[980] = 10'b0001000000;
assign label_2[981] = 10'b0001000000;
assign label_2[982] = 10'b0001000000;
assign label_2[983] = 10'b0001000000;
assign label_2[984] = 10'b0100000000;
assign label_2[985] = 10'b0010000000;
assign label_2[986] = 10'b0100000000;
assign label_2[987] = 10'b0000000100;
assign label_2[988] = 10'b0100000000;
assign label_2[989] = 10'b0100000000;
assign label_2[990] = 10'b0100000000;
assign label_2[991] = 10'b0000000100;
assign label_2[992] = 10'b0000100000;
assign label_2[993] = 10'b0000001000;
assign label_2[994] = 10'b0000000001;
assign label_2[995] = 10'b0000000001;
assign label_2[996] = 10'b0000010000;
assign label_2[997] = 10'b0000000100;
assign label_2[998] = 10'b0000010000;
assign label_2[999] = 10'b0000010000;
assign label_2[1000] = 10'b0000010000;
assign label_2[1001] = 10'b0100000000;
assign label_2[1002] = 10'b0010000000;
assign label_2[1003] = 10'b0010000000;
assign label_2[1004] = 10'b0001000000;
assign label_2[1005] = 10'b0001000000;
assign label_2[1006] = 10'b0001000000;
assign label_2[1007] = 10'b0001000000;
assign label_2[1008] = 10'b0010000000;
assign label_2[1009] = 10'b0000000001;
assign label_2[1010] = 10'b0001000000;
assign label_2[1011] = 10'b0000000001;
assign label_2[1012] = 10'b0000001000;
assign label_2[1013] = 10'b0000001000;
assign label_2[1014] = 10'b0000100000;
assign label_2[1015] = 10'b0000000001;
assign label_2[1016] = 10'b0001000000;
assign label_2[1017] = 10'b0100000000;
assign label_2[1018] = 10'b0100000000;
assign label_2[1019] = 10'b0100000000;
assign label_2[1020] = 10'b0000001000;
assign label_2[1021] = 10'b0000001000;
assign label_2[1022] = 10'b0000000100;
assign label_2[1023] = 10'b0001000000;
assign label_3[0] = 10'b0010000000;
assign label_3[1] = 10'b0010000000;
assign label_3[2] = 10'b0000001000;
assign label_3[3] = 10'b1000000000;
assign label_3[4] = 10'b0010000000;
assign label_3[5] = 10'b0000100000;
assign label_3[6] = 10'b1000000000;
assign label_3[7] = 10'b1000000000;
assign label_3[8] = 10'b0000100000;
assign label_3[9] = 10'b0000010000;
assign label_3[10] = 10'b0001000000;
assign label_3[11] = 10'b0000100000;
assign label_3[12] = 10'b0010000000;
assign label_3[13] = 10'b0000010000;
assign label_3[14] = 10'b0000000001;
assign label_3[15] = 10'b0000010000;
assign label_3[16] = 10'b0000000001;
assign label_3[17] = 10'b0000000001;
assign label_3[18] = 10'b0000100000;
assign label_3[19] = 10'b0000001000;
assign label_3[20] = 10'b0000010000;
assign label_3[21] = 10'b1000000000;
assign label_3[22] = 10'b0001000000;
assign label_3[23] = 10'b0000000001;
assign label_3[24] = 10'b0010000000;
assign label_3[25] = 10'b0001000000;
assign label_3[26] = 10'b0000000001;
assign label_3[27] = 10'b0001000000;
assign label_3[28] = 10'b0001000000;
assign label_3[29] = 10'b0000000001;
assign label_3[30] = 10'b0000000001;
assign label_3[31] = 10'b0000000001;
assign label_3[32] = 10'b0000010000;
assign label_3[33] = 10'b0001000000;
assign label_3[34] = 10'b0000100000;
assign label_3[35] = 10'b1000000000;
assign label_3[36] = 10'b0001000000;
assign label_3[37] = 10'b0000100000;
assign label_3[38] = 10'b0000010000;
assign label_3[39] = 10'b0000000100;
assign label_3[40] = 10'b1000000000;
assign label_3[41] = 10'b0000100000;
assign label_3[42] = 10'b0000100000;
assign label_3[43] = 10'b0000100000;
assign label_3[44] = 10'b0000100000;
assign label_3[45] = 10'b0000100000;
assign label_3[46] = 10'b0000100000;
assign label_3[47] = 10'b0100000000;
assign label_3[48] = 10'b0000100000;
assign label_3[49] = 10'b0001000000;
assign label_3[50] = 10'b0000000100;
assign label_3[51] = 10'b0000001000;
assign label_3[52] = 10'b0100000000;
assign label_3[53] = 10'b1000000000;
assign label_3[54] = 10'b0000000001;
assign label_3[55] = 10'b0001000000;
assign label_3[56] = 10'b0001000000;
assign label_3[57] = 10'b0000100000;
assign label_3[58] = 10'b0001000000;
assign label_3[59] = 10'b0000000100;
assign label_3[60] = 10'b0000000001;
assign label_3[61] = 10'b0000000001;
assign label_3[62] = 10'b0100000000;
assign label_3[63] = 10'b0100000000;
assign label_3[64] = 10'b0000100000;
assign label_3[65] = 10'b0000100000;
assign label_3[66] = 10'b0000000010;
assign label_3[67] = 10'b0000000001;
assign label_3[68] = 10'b0000100000;
assign label_3[69] = 10'b0000000100;
assign label_3[70] = 10'b0000001000;
assign label_3[71] = 10'b0000100000;
assign label_3[72] = 10'b0000000010;
assign label_3[73] = 10'b0000000010;
assign label_3[74] = 10'b0000000010;
assign label_3[75] = 10'b0000000010;
assign label_3[76] = 10'b0000000100;
assign label_3[77] = 10'b0000000100;
assign label_3[78] = 10'b0000000100;
assign label_3[79] = 10'b0000000100;
assign label_3[80] = 10'b0000000001;
assign label_3[81] = 10'b0000000100;
assign label_3[82] = 10'b0000000100;
assign label_3[83] = 10'b0000000100;
assign label_3[84] = 10'b0000010000;
assign label_3[85] = 10'b0000100000;
assign label_3[86] = 10'b0000000100;
assign label_3[87] = 10'b0000000100;
assign label_3[88] = 10'b0000000001;
assign label_3[89] = 10'b0000100000;
assign label_3[90] = 10'b0000000001;
assign label_3[91] = 10'b0000001000;
assign label_3[92] = 10'b0000000001;
assign label_3[93] = 10'b0000000001;
assign label_3[94] = 10'b0000000001;
assign label_3[95] = 10'b0000000001;
assign label_3[96] = 10'b0000001000;
assign label_3[97] = 10'b0000001000;
assign label_3[98] = 10'b0000000001;
assign label_3[99] = 10'b0000001000;
assign label_3[100] = 10'b0000000100;
assign label_3[101] = 10'b0000000001;
assign label_3[102] = 10'b0001000000;
assign label_3[103] = 10'b0000000001;
assign label_3[104] = 10'b0000000001;
assign label_3[105] = 10'b0000010000;
assign label_3[106] = 10'b0000000100;
assign label_3[107] = 10'b0000000100;
assign label_3[108] = 10'b0000100000;
assign label_3[109] = 10'b0000001000;
assign label_3[110] = 10'b0000001000;
assign label_3[111] = 10'b0000001000;
assign label_3[112] = 10'b0000100000;
assign label_3[113] = 10'b0000000100;
assign label_3[114] = 10'b0001000000;
assign label_3[115] = 10'b0000000001;
assign label_3[116] = 10'b0000001000;
assign label_3[117] = 10'b0000100000;
assign label_3[118] = 10'b0000000001;
assign label_3[119] = 10'b0000100000;
assign label_3[120] = 10'b0000100000;
assign label_3[121] = 10'b0000000001;
assign label_3[122] = 10'b0000000001;
assign label_3[123] = 10'b0000000001;
assign label_3[124] = 10'b0000001000;
assign label_3[125] = 10'b0000100000;
assign label_3[126] = 10'b0000000001;
assign label_3[127] = 10'b0000100000;
assign label_3[128] = 10'b0000000010;
assign label_3[129] = 10'b0000010000;
assign label_3[130] = 10'b0000100000;
assign label_3[131] = 10'b0001000000;
assign label_3[132] = 10'b0001000000;
assign label_3[133] = 10'b0010000000;
assign label_3[134] = 10'b0100000000;
assign label_3[135] = 10'b0001000000;
assign label_3[136] = 10'b0000000010;
assign label_3[137] = 10'b0000000100;
assign label_3[138] = 10'b0010000000;
assign label_3[139] = 10'b0000000100;
assign label_3[140] = 10'b1000000000;
assign label_3[141] = 10'b0001000000;
assign label_3[142] = 10'b0001000000;
assign label_3[143] = 10'b0001000000;
assign label_3[144] = 10'b0000000010;
assign label_3[145] = 10'b0000000100;
assign label_3[146] = 10'b0010000000;
assign label_3[147] = 10'b0000000100;
assign label_3[148] = 10'b1000000000;
assign label_3[149] = 10'b0010000000;
assign label_3[150] = 10'b0001000000;
assign label_3[151] = 10'b1000000000;
assign label_3[152] = 10'b0100000000;
assign label_3[153] = 10'b0100000000;
assign label_3[154] = 10'b0010000000;
assign label_3[155] = 10'b0100000000;
assign label_3[156] = 10'b0000000001;
assign label_3[157] = 10'b0000100000;
assign label_3[158] = 10'b0000001000;
assign label_3[159] = 10'b0100000000;
assign label_3[160] = 10'b0000010000;
assign label_3[161] = 10'b0000001000;
assign label_3[162] = 10'b0000010000;
assign label_3[163] = 10'b0001000000;
assign label_3[164] = 10'b1000000000;
assign label_3[165] = 10'b0000100000;
assign label_3[166] = 10'b0000001000;
assign label_3[167] = 10'b0000100000;
assign label_3[168] = 10'b0000001000;
assign label_3[169] = 10'b0000100000;
assign label_3[170] = 10'b0100000000;
assign label_3[171] = 10'b0001000000;
assign label_3[172] = 10'b0000100000;
assign label_3[173] = 10'b0000001000;
assign label_3[174] = 10'b0000100000;
assign label_3[175] = 10'b0100000000;
assign label_3[176] = 10'b0100000000;
assign label_3[177] = 10'b0001000000;
assign label_3[178] = 10'b0001000000;
assign label_3[179] = 10'b0100000000;
assign label_3[180] = 10'b0100000000;
assign label_3[181] = 10'b0000100000;
assign label_3[182] = 10'b0001000000;
assign label_3[183] = 10'b0001000000;
assign label_3[184] = 10'b0100000000;
assign label_3[185] = 10'b0100000000;
assign label_3[186] = 10'b0001000000;
assign label_3[187] = 10'b0100000000;
assign label_3[188] = 10'b0001000000;
assign label_3[189] = 10'b0100000000;
assign label_3[190] = 10'b0001000000;
assign label_3[191] = 10'b0000001000;
assign label_3[192] = 10'b0010000000;
assign label_3[193] = 10'b1000000000;
assign label_3[194] = 10'b0100000000;
assign label_3[195] = 10'b0000000010;
assign label_3[196] = 10'b1000000000;
assign label_3[197] = 10'b0000001000;
assign label_3[198] = 10'b0000000010;
assign label_3[199] = 10'b0100000000;
assign label_3[200] = 10'b0000010000;
assign label_3[201] = 10'b0010000000;
assign label_3[202] = 10'b1000000000;
assign label_3[203] = 10'b0000010000;
assign label_3[204] = 10'b0000000100;
assign label_3[205] = 10'b0010000000;
assign label_3[206] = 10'b0000010000;
assign label_3[207] = 10'b0001000000;
assign label_3[208] = 10'b0000010000;
assign label_3[209] = 10'b0000010000;
assign label_3[210] = 10'b1000000000;
assign label_3[211] = 10'b0000010000;
assign label_3[212] = 10'b0000100000;
assign label_3[213] = 10'b0000010000;
assign label_3[214] = 10'b0000010000;
assign label_3[215] = 10'b1000000000;
assign label_3[216] = 10'b1000000000;
assign label_3[217] = 10'b0001000000;
assign label_3[218] = 10'b0000100000;
assign label_3[219] = 10'b0000001000;
assign label_3[220] = 10'b1000000000;
assign label_3[221] = 10'b0000010000;
assign label_3[222] = 10'b1000000000;
assign label_3[223] = 10'b0100000000;
assign label_3[224] = 10'b0000100000;
assign label_3[225] = 10'b0001000000;
assign label_3[226] = 10'b0000100000;
assign label_3[227] = 10'b0000100000;
assign label_3[228] = 10'b0001000000;
assign label_3[229] = 10'b0000100000;
assign label_3[230] = 10'b0001000000;
assign label_3[231] = 10'b0000000100;
assign label_3[232] = 10'b0000100000;
assign label_3[233] = 10'b0000000001;
assign label_3[234] = 10'b0001000000;
assign label_3[235] = 10'b0000100000;
assign label_3[236] = 10'b0000001000;
assign label_3[237] = 10'b0000100000;
assign label_3[238] = 10'b0000000001;
assign label_3[239] = 10'b0000000001;
assign label_3[240] = 10'b0000100000;
assign label_3[241] = 10'b0000000100;
assign label_3[242] = 10'b0100000000;
assign label_3[243] = 10'b0000000100;
assign label_3[244] = 10'b0000100000;
assign label_3[245] = 10'b0000001000;
assign label_3[246] = 10'b0000100000;
assign label_3[247] = 10'b0100000000;
assign label_3[248] = 10'b0000000100;
assign label_3[249] = 10'b0000010000;
assign label_3[250] = 10'b0000010000;
assign label_3[251] = 10'b0000000100;
assign label_3[252] = 10'b0001000000;
assign label_3[253] = 10'b0000000100;
assign label_3[254] = 10'b1000000000;
assign label_3[255] = 10'b0100000000;
assign label_3[256] = 10'b0010000000;
assign label_3[257] = 10'b0010000000;
assign label_3[258] = 10'b0010000000;
assign label_3[259] = 10'b0010000000;
assign label_3[260] = 10'b0010000000;
assign label_3[261] = 10'b0010000000;
assign label_3[262] = 10'b0010000000;
assign label_3[263] = 10'b0010000000;
assign label_3[264] = 10'b0010000000;
assign label_3[265] = 10'b0010000000;
assign label_3[266] = 10'b0010000000;
assign label_3[267] = 10'b0010000000;
assign label_3[268] = 10'b0010000000;
assign label_3[269] = 10'b0010000000;
assign label_3[270] = 10'b0010000000;
assign label_3[271] = 10'b0010000000;
assign label_3[272] = 10'b0010000000;
assign label_3[273] = 10'b0010000000;
assign label_3[274] = 10'b0010000000;
assign label_3[275] = 10'b0010000000;
assign label_3[276] = 10'b0010000000;
assign label_3[277] = 10'b0010000000;
assign label_3[278] = 10'b0010000000;
assign label_3[279] = 10'b0010000000;
assign label_3[280] = 10'b1000000000;
assign label_3[281] = 10'b1000000000;
assign label_3[282] = 10'b1000000000;
assign label_3[283] = 10'b1000000000;
assign label_3[284] = 10'b1000000000;
assign label_3[285] = 10'b1000000000;
assign label_3[286] = 10'b1000000000;
assign label_3[287] = 10'b1000000000;
assign label_3[288] = 10'b0010000000;
assign label_3[289] = 10'b0010000000;
assign label_3[290] = 10'b1000000000;
assign label_3[291] = 10'b0010000000;
assign label_3[292] = 10'b0010000000;
assign label_3[293] = 10'b0010000000;
assign label_3[294] = 10'b0010000000;
assign label_3[295] = 10'b0010000000;
assign label_3[296] = 10'b1000000000;
assign label_3[297] = 10'b1000000000;
assign label_3[298] = 10'b1000000000;
assign label_3[299] = 10'b1000000000;
assign label_3[300] = 10'b0010000000;
assign label_3[301] = 10'b0010000000;
assign label_3[302] = 10'b0010000000;
assign label_3[303] = 10'b0010000000;
assign label_3[304] = 10'b1000000000;
assign label_3[305] = 10'b0010000000;
assign label_3[306] = 10'b0010000000;
assign label_3[307] = 10'b0010000000;
assign label_3[308] = 10'b1000000000;
assign label_3[309] = 10'b1000000000;
assign label_3[310] = 10'b1000000000;
assign label_3[311] = 10'b1000000000;
assign label_3[312] = 10'b0010000000;
assign label_3[313] = 10'b0010000000;
assign label_3[314] = 10'b0010000000;
assign label_3[315] = 10'b0010000000;
assign label_3[316] = 10'b0010000000;
assign label_3[317] = 10'b0010000000;
assign label_3[318] = 10'b1000000000;
assign label_3[319] = 10'b1000000000;
assign label_3[320] = 10'b0000100000;
assign label_3[321] = 10'b0000100000;
assign label_3[322] = 10'b0000100000;
assign label_3[323] = 10'b0000100000;
assign label_3[324] = 10'b0000100000;
assign label_3[325] = 10'b0000100000;
assign label_3[326] = 10'b0000100000;
assign label_3[327] = 10'b0000100000;
assign label_3[328] = 10'b0010000000;
assign label_3[329] = 10'b0010000000;
assign label_3[330] = 10'b0010000000;
assign label_3[331] = 10'b0010000000;
assign label_3[332] = 10'b0010000000;
assign label_3[333] = 10'b1000000000;
assign label_3[334] = 10'b0010000000;
assign label_3[335] = 10'b0010000000;
assign label_3[336] = 10'b1000000000;
assign label_3[337] = 10'b1000000000;
assign label_3[338] = 10'b1000000000;
assign label_3[339] = 10'b1000000000;
assign label_3[340] = 10'b1000000000;
assign label_3[341] = 10'b1000000000;
assign label_3[342] = 10'b1000000000;
assign label_3[343] = 10'b1000000000;
assign label_3[344] = 10'b0000001000;
assign label_3[345] = 10'b0000001000;
assign label_3[346] = 10'b0000001000;
assign label_3[347] = 10'b0000001000;
assign label_3[348] = 10'b1000000000;
assign label_3[349] = 10'b1000000000;
assign label_3[350] = 10'b1000000000;
assign label_3[351] = 10'b1000000000;
assign label_3[352] = 10'b0010000000;
assign label_3[353] = 10'b0010000000;
assign label_3[354] = 10'b0010000000;
assign label_3[355] = 10'b0010000000;
assign label_3[356] = 10'b0010000000;
assign label_3[357] = 10'b1000000000;
assign label_3[358] = 10'b1000000000;
assign label_3[359] = 10'b1000000000;
assign label_3[360] = 10'b0000100000;
assign label_3[361] = 10'b0000100000;
assign label_3[362] = 10'b0000100000;
assign label_3[363] = 10'b0000100000;
assign label_3[364] = 10'b1000000000;
assign label_3[365] = 10'b0010000000;
assign label_3[366] = 10'b1000000000;
assign label_3[367] = 10'b1000000000;
assign label_3[368] = 10'b0010000000;
assign label_3[369] = 10'b0010000000;
assign label_3[370] = 10'b0010000000;
assign label_3[371] = 10'b0010000000;
assign label_3[372] = 10'b0010000000;
assign label_3[373] = 10'b0010000000;
assign label_3[374] = 10'b0010000000;
assign label_3[375] = 10'b0010000000;
assign label_3[376] = 10'b1000000000;
assign label_3[377] = 10'b1000000000;
assign label_3[378] = 10'b0010000000;
assign label_3[379] = 10'b0010000000;
assign label_3[380] = 10'b0010000000;
assign label_3[381] = 10'b0100000000;
assign label_3[382] = 10'b1000000000;
assign label_3[383] = 10'b1000000000;
assign label_3[384] = 10'b0010000000;
assign label_3[385] = 10'b0010000000;
assign label_3[386] = 10'b0010000000;
assign label_3[387] = 10'b1000000000;
assign label_3[388] = 10'b0010000000;
assign label_3[389] = 10'b0010000000;
assign label_3[390] = 10'b0000010000;
assign label_3[391] = 10'b0010000000;
assign label_3[392] = 10'b0000100000;
assign label_3[393] = 10'b0000100000;
assign label_3[394] = 10'b0000100000;
assign label_3[395] = 10'b0000100000;
assign label_3[396] = 10'b0000100000;
assign label_3[397] = 10'b0000100000;
assign label_3[398] = 10'b0000100000;
assign label_3[399] = 10'b0000100000;
assign label_3[400] = 10'b0010000000;
assign label_3[401] = 10'b0010000000;
assign label_3[402] = 10'b0000001000;
assign label_3[403] = 10'b1000000000;
assign label_3[404] = 10'b0010000000;
assign label_3[405] = 10'b0010000000;
assign label_3[406] = 10'b0010000000;
assign label_3[407] = 10'b0010000000;
assign label_3[408] = 10'b0010000000;
assign label_3[409] = 10'b0010000000;
assign label_3[410] = 10'b1000000000;
assign label_3[411] = 10'b1000000000;
assign label_3[412] = 10'b0010000000;
assign label_3[413] = 10'b0010000000;
assign label_3[414] = 10'b1000000000;
assign label_3[415] = 10'b0010000000;
assign label_3[416] = 10'b1000000000;
assign label_3[417] = 10'b1000000000;
assign label_3[418] = 10'b1000000000;
assign label_3[419] = 10'b1000000000;
assign label_3[420] = 10'b1000000000;
assign label_3[421] = 10'b1000000000;
assign label_3[422] = 10'b1000000000;
assign label_3[423] = 10'b1000000000;
assign label_3[424] = 10'b0010000000;
assign label_3[425] = 10'b0010000000;
assign label_3[426] = 10'b0010000000;
assign label_3[427] = 10'b0010000000;
assign label_3[428] = 10'b1000000000;
assign label_3[429] = 10'b0010000000;
assign label_3[430] = 10'b1000000000;
assign label_3[431] = 10'b1000000000;
assign label_3[432] = 10'b0000001000;
assign label_3[433] = 10'b0000001000;
assign label_3[434] = 10'b0000001000;
assign label_3[435] = 10'b0000001000;
assign label_3[436] = 10'b0010000000;
assign label_3[437] = 10'b0010000000;
assign label_3[438] = 10'b0010000000;
assign label_3[439] = 10'b0010000000;
assign label_3[440] = 10'b0000100000;
assign label_3[441] = 10'b0000100000;
assign label_3[442] = 10'b0000100000;
assign label_3[443] = 10'b0000100000;
assign label_3[444] = 10'b1000000000;
assign label_3[445] = 10'b0100000000;
assign label_3[446] = 10'b0010000000;
assign label_3[447] = 10'b0010000000;
assign label_3[448] = 10'b1000000000;
assign label_3[449] = 10'b1000000000;
assign label_3[450] = 10'b1000000000;
assign label_3[451] = 10'b1000000000;
assign label_3[452] = 10'b0000100000;
assign label_3[453] = 10'b0000100000;
assign label_3[454] = 10'b0000100000;
assign label_3[455] = 10'b0000100000;
assign label_3[456] = 10'b1000000000;
assign label_3[457] = 10'b1000000000;
assign label_3[458] = 10'b1000000000;
assign label_3[459] = 10'b1000000000;
assign label_3[460] = 10'b0000100000;
assign label_3[461] = 10'b0000100000;
assign label_3[462] = 10'b0000100000;
assign label_3[463] = 10'b0000100000;
assign label_3[464] = 10'b0010000000;
assign label_3[465] = 10'b0010000000;
assign label_3[466] = 10'b0010000000;
assign label_3[467] = 10'b0010000000;
assign label_3[468] = 10'b0000010000;
assign label_3[469] = 10'b1000000000;
assign label_3[470] = 10'b0010000000;
assign label_3[471] = 10'b0010000000;
assign label_3[472] = 10'b0100000000;
assign label_3[473] = 10'b1000000000;
assign label_3[474] = 10'b1000000000;
assign label_3[475] = 10'b1000000000;
assign label_3[476] = 10'b1000000000;
assign label_3[477] = 10'b1000000000;
assign label_3[478] = 10'b0010000000;
assign label_3[479] = 10'b0010000000;
assign label_3[480] = 10'b0010000000;
assign label_3[481] = 10'b0010000000;
assign label_3[482] = 10'b0010000000;
assign label_3[483] = 10'b0010000000;
assign label_3[484] = 10'b0010000000;
assign label_3[485] = 10'b0010000000;
assign label_3[486] = 10'b0010000000;
assign label_3[487] = 10'b0010000000;
assign label_3[488] = 10'b0000100000;
assign label_3[489] = 10'b0000100000;
assign label_3[490] = 10'b0010000000;
assign label_3[491] = 10'b0010000000;
assign label_3[492] = 10'b0000100000;
assign label_3[493] = 10'b0000100000;
assign label_3[494] = 10'b1000000000;
assign label_3[495] = 10'b1000000000;
assign label_3[496] = 10'b1000000000;
assign label_3[497] = 10'b1000000000;
assign label_3[498] = 10'b0000100000;
assign label_3[499] = 10'b0000100000;
assign label_3[500] = 10'b1000000000;
assign label_3[501] = 10'b1000000000;
assign label_3[502] = 10'b1000000000;
assign label_3[503] = 10'b1000000000;
assign label_3[504] = 10'b0000100000;
assign label_3[505] = 10'b0000100000;
assign label_3[506] = 10'b0000100000;
assign label_3[507] = 10'b0000100000;
assign label_3[508] = 10'b0000100000;
assign label_3[509] = 10'b0000100000;
assign label_3[510] = 10'b0000100000;
assign label_3[511] = 10'b0000100000;
assign label_3[512] = 10'b0000001000;
assign label_3[513] = 10'b0000100000;
assign label_3[514] = 10'b0000100000;
assign label_3[515] = 10'b0000100000;
assign label_3[516] = 10'b0000000010;
assign label_3[517] = 10'b0001000000;
assign label_3[518] = 10'b0000000010;
assign label_3[519] = 10'b0000000100;
assign label_3[520] = 10'b0100000000;
assign label_3[521] = 10'b0000000100;
assign label_3[522] = 10'b0000010000;
assign label_3[523] = 10'b0000010000;
assign label_3[524] = 10'b0000100000;
assign label_3[525] = 10'b0000000001;
assign label_3[526] = 10'b0000010000;
assign label_3[527] = 10'b0000100000;
assign label_3[528] = 10'b0000010000;
assign label_3[529] = 10'b0001000000;
assign label_3[530] = 10'b0000100000;
assign label_3[531] = 10'b0000100000;
assign label_3[532] = 10'b0000010000;
assign label_3[533] = 10'b0100000000;
assign label_3[534] = 10'b0000010000;
assign label_3[535] = 10'b1000000000;
assign label_3[536] = 10'b0000000100;
assign label_3[537] = 10'b0000100000;
assign label_3[538] = 10'b0001000000;
assign label_3[539] = 10'b0001000000;
assign label_3[540] = 10'b0000000100;
assign label_3[541] = 10'b0000100000;
assign label_3[542] = 10'b0000000100;
assign label_3[543] = 10'b0000001000;
assign label_3[544] = 10'b0001000000;
assign label_3[545] = 10'b0000010000;
assign label_3[546] = 10'b0000000100;
assign label_3[547] = 10'b0001000000;
assign label_3[548] = 10'b0000000100;
assign label_3[549] = 10'b0000100000;
assign label_3[550] = 10'b0000010000;
assign label_3[551] = 10'b0000000001;
assign label_3[552] = 10'b0000000001;
assign label_3[553] = 10'b0000000100;
assign label_3[554] = 10'b0001000000;
assign label_3[555] = 10'b0000000100;
assign label_3[556] = 10'b0000000100;
assign label_3[557] = 10'b0000000001;
assign label_3[558] = 10'b0001000000;
assign label_3[559] = 10'b0000010000;
assign label_3[560] = 10'b0000000001;
assign label_3[561] = 10'b0100000000;
assign label_3[562] = 10'b0000000010;
assign label_3[563] = 10'b0001000000;
assign label_3[564] = 10'b0000000100;
assign label_3[565] = 10'b0100000000;
assign label_3[566] = 10'b0000000100;
assign label_3[567] = 10'b0000000001;
assign label_3[568] = 10'b0000000001;
assign label_3[569] = 10'b0000000100;
assign label_3[570] = 10'b0000000001;
assign label_3[571] = 10'b0000100000;
assign label_3[572] = 10'b0000000100;
assign label_3[573] = 10'b0001000000;
assign label_3[574] = 10'b0000000100;
assign label_3[575] = 10'b0000000100;
assign label_3[576] = 10'b0000000100;
assign label_3[577] = 10'b0000001000;
assign label_3[578] = 10'b0000000100;
assign label_3[579] = 10'b0000000100;
assign label_3[580] = 10'b0000000001;
assign label_3[581] = 10'b0000000001;
assign label_3[582] = 10'b0001000000;
assign label_3[583] = 10'b0001000000;
assign label_3[584] = 10'b0001000000;
assign label_3[585] = 10'b0001000000;
assign label_3[586] = 10'b0001000000;
assign label_3[587] = 10'b0001000000;
assign label_3[588] = 10'b0001000000;
assign label_3[589] = 10'b0001000000;
assign label_3[590] = 10'b0001000000;
assign label_3[591] = 10'b0001000000;
assign label_3[592] = 10'b0000100000;
assign label_3[593] = 10'b0000100000;
assign label_3[594] = 10'b0000001000;
assign label_3[595] = 10'b0000001000;
assign label_3[596] = 10'b0000001000;
assign label_3[597] = 10'b0000001000;
assign label_3[598] = 10'b0000100000;
assign label_3[599] = 10'b0001000000;
assign label_3[600] = 10'b0000000100;
assign label_3[601] = 10'b0001000000;
assign label_3[602] = 10'b0000100000;
assign label_3[603] = 10'b0000000001;
assign label_3[604] = 10'b0000000100;
assign label_3[605] = 10'b0000000100;
assign label_3[606] = 10'b0000000100;
assign label_3[607] = 10'b0000000100;
assign label_3[608] = 10'b0000000100;
assign label_3[609] = 10'b0000000100;
assign label_3[610] = 10'b0000000100;
assign label_3[611] = 10'b0001000000;
assign label_3[612] = 10'b0000000100;
assign label_3[613] = 10'b0000000100;
assign label_3[614] = 10'b0000100000;
assign label_3[615] = 10'b0001000000;
assign label_3[616] = 10'b0001000000;
assign label_3[617] = 10'b0001000000;
assign label_3[618] = 10'b0000000100;
assign label_3[619] = 10'b0000000100;
assign label_3[620] = 10'b0000001000;
assign label_3[621] = 10'b0000000100;
assign label_3[622] = 10'b0000000001;
assign label_3[623] = 10'b0000010000;
assign label_3[624] = 10'b0000000100;
assign label_3[625] = 10'b0000000100;
assign label_3[626] = 10'b0000000100;
assign label_3[627] = 10'b0000000100;
assign label_3[628] = 10'b0000000100;
assign label_3[629] = 10'b0100000000;
assign label_3[630] = 10'b0000000100;
assign label_3[631] = 10'b0000000100;
assign label_3[632] = 10'b0100000000;
assign label_3[633] = 10'b0000000100;
assign label_3[634] = 10'b0000001000;
assign label_3[635] = 10'b0000001000;
assign label_3[636] = 10'b0000000100;
assign label_3[637] = 10'b0000000100;
assign label_3[638] = 10'b0000100000;
assign label_3[639] = 10'b0000100000;
assign label_3[640] = 10'b0001000000;
assign label_3[641] = 10'b0000100000;
assign label_3[642] = 10'b0000000001;
assign label_3[643] = 10'b0000100000;
assign label_3[644] = 10'b0000000001;
assign label_3[645] = 10'b0000000100;
assign label_3[646] = 10'b0000001000;
assign label_3[647] = 10'b0000000001;
assign label_3[648] = 10'b0000000001;
assign label_3[649] = 10'b0000000100;
assign label_3[650] = 10'b0000100000;
assign label_3[651] = 10'b0000000001;
assign label_3[652] = 10'b0000100000;
assign label_3[653] = 10'b0000001000;
assign label_3[654] = 10'b0000000001;
assign label_3[655] = 10'b0000000001;
assign label_3[656] = 10'b0000000001;
assign label_3[657] = 10'b0000000001;
assign label_3[658] = 10'b0001000000;
assign label_3[659] = 10'b0001000000;
assign label_3[660] = 10'b0000001000;
assign label_3[661] = 10'b0000000001;
assign label_3[662] = 10'b0000000001;
assign label_3[663] = 10'b0000100000;
assign label_3[664] = 10'b0000000100;
assign label_3[665] = 10'b0001000000;
assign label_3[666] = 10'b0001000000;
assign label_3[667] = 10'b0000000001;
assign label_3[668] = 10'b0100000000;
assign label_3[669] = 10'b0000000001;
assign label_3[670] = 10'b0000001000;
assign label_3[671] = 10'b0000001000;
assign label_3[672] = 10'b0001000000;
assign label_3[673] = 10'b0001000000;
assign label_3[674] = 10'b0000000001;
assign label_3[675] = 10'b0000000001;
assign label_3[676] = 10'b0000000100;
assign label_3[677] = 10'b0000000100;
assign label_3[678] = 10'b0100000000;
assign label_3[679] = 10'b0100000000;
assign label_3[680] = 10'b0100000000;
assign label_3[681] = 10'b0100000000;
assign label_3[682] = 10'b0100000000;
assign label_3[683] = 10'b0100000000;
assign label_3[684] = 10'b0100000000;
assign label_3[685] = 10'b0100000000;
assign label_3[686] = 10'b0100000000;
assign label_3[687] = 10'b0100000000;
assign label_3[688] = 10'b0000000100;
assign label_3[689] = 10'b0000000100;
assign label_3[690] = 10'b0000000100;
assign label_3[691] = 10'b0100000000;
assign label_3[692] = 10'b1000000000;
assign label_3[693] = 10'b0000010000;
assign label_3[694] = 10'b0000001000;
assign label_3[695] = 10'b0000001000;
assign label_3[696] = 10'b0000010000;
assign label_3[697] = 10'b0000010000;
assign label_3[698] = 10'b0000010000;
assign label_3[699] = 10'b0000010000;
assign label_3[700] = 10'b0001000000;
assign label_3[701] = 10'b0100000000;
assign label_3[702] = 10'b0000000001;
assign label_3[703] = 10'b0000000001;
assign label_3[704] = 10'b0000000100;
assign label_3[705] = 10'b0000001000;
assign label_3[706] = 10'b0000010000;
assign label_3[707] = 10'b1000000000;
assign label_3[708] = 10'b0100000000;
assign label_3[709] = 10'b0000000100;
assign label_3[710] = 10'b0000001000;
assign label_3[711] = 10'b0001000000;
assign label_3[712] = 10'b0000010000;
assign label_3[713] = 10'b0001000000;
assign label_3[714] = 10'b0001000000;
assign label_3[715] = 10'b0100000000;
assign label_3[716] = 10'b0100000000;
assign label_3[717] = 10'b0100000000;
assign label_3[718] = 10'b1000000000;
assign label_3[719] = 10'b0000000100;
assign label_3[720] = 10'b0000000100;
assign label_3[721] = 10'b0000001000;
assign label_3[722] = 10'b0000000001;
assign label_3[723] = 10'b0000000100;
assign label_3[724] = 10'b0000000100;
assign label_3[725] = 10'b0001000000;
assign label_3[726] = 10'b1000000000;
assign label_3[727] = 10'b1000000000;
assign label_3[728] = 10'b0100000000;
assign label_3[729] = 10'b0100000000;
assign label_3[730] = 10'b0100000000;
assign label_3[731] = 10'b0100000000;
assign label_3[732] = 10'b0001000000;
assign label_3[733] = 10'b0001000000;
assign label_3[734] = 10'b0001000000;
assign label_3[735] = 10'b0001000000;
assign label_3[736] = 10'b0001000000;
assign label_3[737] = 10'b0000010000;
assign label_3[738] = 10'b0100000000;
assign label_3[739] = 10'b1000000000;
assign label_3[740] = 10'b0001000000;
assign label_3[741] = 10'b0000010000;
assign label_3[742] = 10'b0001000000;
assign label_3[743] = 10'b0000000001;
assign label_3[744] = 10'b0000010000;
assign label_3[745] = 10'b0000010000;
assign label_3[746] = 10'b0000100000;
assign label_3[747] = 10'b0000100000;
assign label_3[748] = 10'b0000001000;
assign label_3[749] = 10'b0000001000;
assign label_3[750] = 10'b1000000000;
assign label_3[751] = 10'b0000000001;
assign label_3[752] = 10'b0000000100;
assign label_3[753] = 10'b0000000100;
assign label_3[754] = 10'b0000000100;
assign label_3[755] = 10'b0000000100;
assign label_3[756] = 10'b1000000000;
assign label_3[757] = 10'b1000000000;
assign label_3[758] = 10'b0100000000;
assign label_3[759] = 10'b0100000000;
assign label_3[760] = 10'b0001000000;
assign label_3[761] = 10'b0001000000;
assign label_3[762] = 10'b0100000000;
assign label_3[763] = 10'b0000000001;
assign label_3[764] = 10'b0000000001;
assign label_3[765] = 10'b0001000000;
assign label_3[766] = 10'b0000000001;
assign label_3[767] = 10'b1000000000;
assign label_3[768] = 10'b0000001000;
assign label_3[769] = 10'b0000000100;
assign label_3[770] = 10'b0000000010;
assign label_3[771] = 10'b0100000000;
assign label_3[772] = 10'b0000000010;
assign label_3[773] = 10'b0000000010;
assign label_3[774] = 10'b0000000100;
assign label_3[775] = 10'b0000001000;
assign label_3[776] = 10'b0000001000;
assign label_3[777] = 10'b0000100000;
assign label_3[778] = 10'b0100000000;
assign label_3[779] = 10'b0100000000;
assign label_3[780] = 10'b0000001000;
assign label_3[781] = 10'b0000000010;
assign label_3[782] = 10'b0000001000;
assign label_3[783] = 10'b0000001000;
assign label_3[784] = 10'b0000000100;
assign label_3[785] = 10'b0000001000;
assign label_3[786] = 10'b0100000000;
assign label_3[787] = 10'b0000100000;
assign label_3[788] = 10'b0100000000;
assign label_3[789] = 10'b0100000000;
assign label_3[790] = 10'b0000000010;
assign label_3[791] = 10'b0000001000;
assign label_3[792] = 10'b0000001000;
assign label_3[793] = 10'b0100000000;
assign label_3[794] = 10'b0000000100;
assign label_3[795] = 10'b0000000100;
assign label_3[796] = 10'b0000001000;
assign label_3[797] = 10'b0100000000;
assign label_3[798] = 10'b0000100000;
assign label_3[799] = 10'b0000100000;
assign label_3[800] = 10'b0000001000;
assign label_3[801] = 10'b0000000010;
assign label_3[802] = 10'b0000001000;
assign label_3[803] = 10'b0000001000;
assign label_3[804] = 10'b0000001000;
assign label_3[805] = 10'b0000001000;
assign label_3[806] = 10'b0000000100;
assign label_3[807] = 10'b0000001000;
assign label_3[808] = 10'b0100000000;
assign label_3[809] = 10'b0000001000;
assign label_3[810] = 10'b0000001000;
assign label_3[811] = 10'b0100000000;
assign label_3[812] = 10'b0001000000;
assign label_3[813] = 10'b0000000100;
assign label_3[814] = 10'b0000001000;
assign label_3[815] = 10'b0000000100;
assign label_3[816] = 10'b0000001000;
assign label_3[817] = 10'b0000100000;
assign label_3[818] = 10'b0000001000;
assign label_3[819] = 10'b0000001000;
assign label_3[820] = 10'b0000100000;
assign label_3[821] = 10'b0000001000;
assign label_3[822] = 10'b0000000001;
assign label_3[823] = 10'b0000000001;
assign label_3[824] = 10'b0100000000;
assign label_3[825] = 10'b0000001000;
assign label_3[826] = 10'b0001000000;
assign label_3[827] = 10'b0001000000;
assign label_3[828] = 10'b0100000000;
assign label_3[829] = 10'b0000000100;
assign label_3[830] = 10'b0000001000;
assign label_3[831] = 10'b0000000001;
assign label_3[832] = 10'b0000000010;
assign label_3[833] = 10'b0000000100;
assign label_3[834] = 10'b0000001000;
assign label_3[835] = 10'b0000000100;
assign label_3[836] = 10'b0100000000;
assign label_3[837] = 10'b0000100000;
assign label_3[838] = 10'b0001000000;
assign label_3[839] = 10'b0000010000;
assign label_3[840] = 10'b0000000100;
assign label_3[841] = 10'b0000000100;
assign label_3[842] = 10'b0000001000;
assign label_3[843] = 10'b0000100000;
assign label_3[844] = 10'b0001000000;
assign label_3[845] = 10'b0001000000;
assign label_3[846] = 10'b0001000000;
assign label_3[847] = 10'b0001000000;
assign label_3[848] = 10'b0001000000;
assign label_3[849] = 10'b0001000000;
assign label_3[850] = 10'b0100000000;
assign label_3[851] = 10'b0100000000;
assign label_3[852] = 10'b0000000100;
assign label_3[853] = 10'b0000010000;
assign label_3[854] = 10'b1000000000;
assign label_3[855] = 10'b0100000000;
assign label_3[856] = 10'b0000010000;
assign label_3[857] = 10'b0000010000;
assign label_3[858] = 10'b0001000000;
assign label_3[859] = 10'b0000000001;
assign label_3[860] = 10'b0100000000;
assign label_3[861] = 10'b0000000100;
assign label_3[862] = 10'b0000001000;
assign label_3[863] = 10'b0000001000;
assign label_3[864] = 10'b0000001000;
assign label_3[865] = 10'b0000001000;
assign label_3[866] = 10'b0100000000;
assign label_3[867] = 10'b0000001000;
assign label_3[868] = 10'b0100000000;
assign label_3[869] = 10'b0000000100;
assign label_3[870] = 10'b0000000100;
assign label_3[871] = 10'b0000000100;
assign label_3[872] = 10'b0100000000;
assign label_3[873] = 10'b0000000010;
assign label_3[874] = 10'b0100000000;
assign label_3[875] = 10'b0100000000;
assign label_3[876] = 10'b0000000100;
assign label_3[877] = 10'b0100000000;
assign label_3[878] = 10'b0100000000;
assign label_3[879] = 10'b0000000100;
assign label_3[880] = 10'b0000001000;
assign label_3[881] = 10'b0000001000;
assign label_3[882] = 10'b0000001000;
assign label_3[883] = 10'b0000001000;
assign label_3[884] = 10'b0000001000;
assign label_3[885] = 10'b0000001000;
assign label_3[886] = 10'b0000000100;
assign label_3[887] = 10'b0000000100;
assign label_3[888] = 10'b0000000100;
assign label_3[889] = 10'b0000000100;
assign label_3[890] = 10'b0000000100;
assign label_3[891] = 10'b0000000100;
assign label_3[892] = 10'b0000000100;
assign label_3[893] = 10'b0000000100;
assign label_3[894] = 10'b0000000100;
assign label_3[895] = 10'b0000000100;
assign label_3[896] = 10'b0000001000;
assign label_3[897] = 10'b0000100000;
assign label_3[898] = 10'b0000001000;
assign label_3[899] = 10'b0100000000;
assign label_3[900] = 10'b0000010000;
assign label_3[901] = 10'b0000100000;
assign label_3[902] = 10'b0100000000;
assign label_3[903] = 10'b0000001000;
assign label_3[904] = 10'b0000000100;
assign label_3[905] = 10'b0000000100;
assign label_3[906] = 10'b0000000100;
assign label_3[907] = 10'b0000000100;
assign label_3[908] = 10'b0000001000;
assign label_3[909] = 10'b0100000000;
assign label_3[910] = 10'b0000001000;
assign label_3[911] = 10'b0000000100;
assign label_3[912] = 10'b0000100000;
assign label_3[913] = 10'b0000001000;
assign label_3[914] = 10'b0000100000;
assign label_3[915] = 10'b0000100000;
assign label_3[916] = 10'b0000001000;
assign label_3[917] = 10'b0000001000;
assign label_3[918] = 10'b0000001000;
assign label_3[919] = 10'b0000000001;
assign label_3[920] = 10'b0001000000;
assign label_3[921] = 10'b0000000001;
assign label_3[922] = 10'b0000000001;
assign label_3[923] = 10'b0001000000;
assign label_3[924] = 10'b0000010000;
assign label_3[925] = 10'b0100000000;
assign label_3[926] = 10'b0001000000;
assign label_3[927] = 10'b0000001000;
assign label_3[928] = 10'b0000100000;
assign label_3[929] = 10'b0001000000;
assign label_3[930] = 10'b0100000000;
assign label_3[931] = 10'b0000001000;
assign label_3[932] = 10'b0000100000;
assign label_3[933] = 10'b0000100000;
assign label_3[934] = 10'b0001000000;
assign label_3[935] = 10'b0000100000;
assign label_3[936] = 10'b0000100000;
assign label_3[937] = 10'b0000100000;
assign label_3[938] = 10'b0100000000;
assign label_3[939] = 10'b0000100000;
assign label_3[940] = 10'b0100000000;
assign label_3[941] = 10'b0000001000;
assign label_3[942] = 10'b0000100000;
assign label_3[943] = 10'b0100000000;
assign label_3[944] = 10'b0000100000;
assign label_3[945] = 10'b0100000000;
assign label_3[946] = 10'b0100000000;
assign label_3[947] = 10'b0000001000;
assign label_3[948] = 10'b0000010000;
assign label_3[949] = 10'b0000010000;
assign label_3[950] = 10'b0100000000;
assign label_3[951] = 10'b0000000001;
assign label_3[952] = 10'b0000100000;
assign label_3[953] = 10'b0000100000;
assign label_3[954] = 10'b0000100000;
assign label_3[955] = 10'b0000100000;
assign label_3[956] = 10'b0000100000;
assign label_3[957] = 10'b0001000000;
assign label_3[958] = 10'b0000000001;
assign label_3[959] = 10'b0000000001;
assign label_3[960] = 10'b0000000100;
assign label_3[961] = 10'b0000100000;
assign label_3[962] = 10'b0000100000;
assign label_3[963] = 10'b0000010000;
assign label_3[964] = 10'b0000001000;
assign label_3[965] = 10'b0000001000;
assign label_3[966] = 10'b0000001000;
assign label_3[967] = 10'b0000001000;
assign label_3[968] = 10'b0000001000;
assign label_3[969] = 10'b0000000100;
assign label_3[970] = 10'b0000001000;
assign label_3[971] = 10'b0100000000;
assign label_3[972] = 10'b0001000000;
assign label_3[973] = 10'b0100000000;
assign label_3[974] = 10'b0000000001;
assign label_3[975] = 10'b0100000000;
assign label_3[976] = 10'b0001000000;
assign label_3[977] = 10'b0100000000;
assign label_3[978] = 10'b0001000000;
assign label_3[979] = 10'b0000000100;
assign label_3[980] = 10'b0100000000;
assign label_3[981] = 10'b0000000010;
assign label_3[982] = 10'b0100000000;
assign label_3[983] = 10'b0100000000;
assign label_3[984] = 10'b0001000000;
assign label_3[985] = 10'b0100000000;
assign label_3[986] = 10'b0100000000;
assign label_3[987] = 10'b0000000001;
assign label_3[988] = 10'b0000000100;
assign label_3[989] = 10'b0100000000;
assign label_3[990] = 10'b0000000001;
assign label_3[991] = 10'b0100000000;
assign label_3[992] = 10'b0100000000;
assign label_3[993] = 10'b0100000000;
assign label_3[994] = 10'b0000100000;
assign label_3[995] = 10'b0000001000;
assign label_3[996] = 10'b0000001000;
assign label_3[997] = 10'b0000100000;
assign label_3[998] = 10'b1000000000;
assign label_3[999] = 10'b1000000000;
assign label_3[1000] = 10'b0100000000;
assign label_3[1001] = 10'b0000001000;
assign label_3[1002] = 10'b0001000000;
assign label_3[1003] = 10'b0000001000;
assign label_3[1004] = 10'b0100000000;
assign label_3[1005] = 10'b0001000000;
assign label_3[1006] = 10'b0000000100;
assign label_3[1007] = 10'b0000000100;
assign label_3[1008] = 10'b1000000000;
assign label_3[1009] = 10'b0000100000;
assign label_3[1010] = 10'b0001000000;
assign label_3[1011] = 10'b0000000100;
assign label_3[1012] = 10'b0000001000;
assign label_3[1013] = 10'b0100000000;
assign label_3[1014] = 10'b0000000001;
assign label_3[1015] = 10'b0100000000;
assign label_3[1016] = 10'b0000100000;
assign label_3[1017] = 10'b0001000000;
assign label_3[1018] = 10'b0001000000;
assign label_3[1019] = 10'b0100000000;
assign label_3[1020] = 10'b0100000000;
assign label_3[1021] = 10'b0000010000;
assign label_3[1022] = 10'b0001000000;
assign label_3[1023] = 10'b0000000001;
assign label_4[0] = 10'b0000000010;
assign label_4[1] = 10'b0000000100;
assign label_4[2] = 10'b0000001000;
assign label_4[3] = 10'b0000000010;
assign label_4[4] = 10'b0000000100;
assign label_4[5] = 10'b0000001000;
assign label_4[6] = 10'b0010000000;
assign label_4[7] = 10'b0001000000;
assign label_4[8] = 10'b0000100000;
assign label_4[9] = 10'b0001000000;
assign label_4[10] = 10'b0000000001;
assign label_4[11] = 10'b0000000001;
assign label_4[12] = 10'b0100000000;
assign label_4[13] = 10'b0000000010;
assign label_4[14] = 10'b0000100000;
assign label_4[15] = 10'b0100000000;
assign label_4[16] = 10'b0001000000;
assign label_4[17] = 10'b0010000000;
assign label_4[18] = 10'b0000000001;
assign label_4[19] = 10'b0000001000;
assign label_4[20] = 10'b0010000000;
assign label_4[21] = 10'b0010000000;
assign label_4[22] = 10'b0010000000;
assign label_4[23] = 10'b0010000000;
assign label_4[24] = 10'b0000000100;
assign label_4[25] = 10'b0001000000;
assign label_4[26] = 10'b0000010000;
assign label_4[27] = 10'b0000000100;
assign label_4[28] = 10'b0000010000;
assign label_4[29] = 10'b0000000100;
assign label_4[30] = 10'b0000001000;
assign label_4[31] = 10'b0000001000;
assign label_4[32] = 10'b0000100000;
assign label_4[33] = 10'b0000001000;
assign label_4[34] = 10'b0000100000;
assign label_4[35] = 10'b0000000001;
assign label_4[36] = 10'b0000000010;
assign label_4[37] = 10'b0000000010;
assign label_4[38] = 10'b0001000000;
assign label_4[39] = 10'b0001000000;
assign label_4[40] = 10'b0000100000;
assign label_4[41] = 10'b0000000001;
assign label_4[42] = 10'b0010000000;
assign label_4[43] = 10'b0000001000;
assign label_4[44] = 10'b0010000000;
assign label_4[45] = 10'b0000000001;
assign label_4[46] = 10'b0000000100;
assign label_4[47] = 10'b0000000100;
assign label_4[48] = 10'b0000100000;
assign label_4[49] = 10'b0000001000;
assign label_4[50] = 10'b0010000000;
assign label_4[51] = 10'b0000100000;
assign label_4[52] = 10'b0000010000;
assign label_4[53] = 10'b1000000000;
assign label_4[54] = 10'b0000000010;
assign label_4[55] = 10'b0010000000;
assign label_4[56] = 10'b1000000000;
assign label_4[57] = 10'b0100000000;
assign label_4[58] = 10'b0100000000;
assign label_4[59] = 10'b0100000000;
assign label_4[60] = 10'b0100000000;
assign label_4[61] = 10'b0100000000;
assign label_4[62] = 10'b0000001000;
assign label_4[63] = 10'b0100000000;
assign label_4[64] = 10'b0010000000;
assign label_4[65] = 10'b0000000100;
assign label_4[66] = 10'b0000010000;
assign label_4[67] = 10'b1000000000;
assign label_4[68] = 10'b0000000100;
assign label_4[69] = 10'b0000001000;
assign label_4[70] = 10'b0000000001;
assign label_4[71] = 10'b0001000000;
assign label_4[72] = 10'b0010000000;
assign label_4[73] = 10'b0000001000;
assign label_4[74] = 10'b0000000010;
assign label_4[75] = 10'b0000100000;
assign label_4[76] = 10'b0010000000;
assign label_4[77] = 10'b0000000100;
assign label_4[78] = 10'b0100000000;
assign label_4[79] = 10'b0100000000;
assign label_4[80] = 10'b0010000000;
assign label_4[81] = 10'b0000000100;
assign label_4[82] = 10'b1000000000;
assign label_4[83] = 10'b0000010000;
assign label_4[84] = 10'b0000000100;
assign label_4[85] = 10'b0000000100;
assign label_4[86] = 10'b0000000100;
assign label_4[87] = 10'b0000000100;
assign label_4[88] = 10'b0000001000;
assign label_4[89] = 10'b0001000000;
assign label_4[90] = 10'b0100000000;
assign label_4[91] = 10'b0000100000;
assign label_4[92] = 10'b0000000100;
assign label_4[93] = 10'b0000000100;
assign label_4[94] = 10'b0001000000;
assign label_4[95] = 10'b0000000100;
assign label_4[96] = 10'b0000001000;
assign label_4[97] = 10'b0000000100;
assign label_4[98] = 10'b0000000100;
assign label_4[99] = 10'b0001000000;
assign label_4[100] = 10'b0000000001;
assign label_4[101] = 10'b0010000000;
assign label_4[102] = 10'b0001000000;
assign label_4[103] = 10'b0000000100;
assign label_4[104] = 10'b0000000100;
assign label_4[105] = 10'b0000010000;
assign label_4[106] = 10'b0000010000;
assign label_4[107] = 10'b0000000100;
assign label_4[108] = 10'b0000000100;
assign label_4[109] = 10'b0001000000;
assign label_4[110] = 10'b0010000000;
assign label_4[111] = 10'b0000000100;
assign label_4[112] = 10'b0000010000;
assign label_4[113] = 10'b0000000001;
assign label_4[114] = 10'b0000000001;
assign label_4[115] = 10'b1000000000;
assign label_4[116] = 10'b1000000000;
assign label_4[117] = 10'b1000000000;
assign label_4[118] = 10'b1000000000;
assign label_4[119] = 10'b1000000000;
assign label_4[120] = 10'b0000000001;
assign label_4[121] = 10'b0000000001;
assign label_4[122] = 10'b0000000001;
assign label_4[123] = 10'b0000000001;
assign label_4[124] = 10'b0001000000;
assign label_4[125] = 10'b0000000001;
assign label_4[126] = 10'b0000000001;
assign label_4[127] = 10'b1000000000;
assign label_4[128] = 10'b0001000000;
assign label_4[129] = 10'b0000010000;
assign label_4[130] = 10'b0000010000;
assign label_4[131] = 10'b0010000000;
assign label_4[132] = 10'b0000000010;
assign label_4[133] = 10'b0000001000;
assign label_4[134] = 10'b0000000100;
assign label_4[135] = 10'b0010000000;
assign label_4[136] = 10'b0000010000;
assign label_4[137] = 10'b0001000000;
assign label_4[138] = 10'b0000010000;
assign label_4[139] = 10'b0000010000;
assign label_4[140] = 10'b0000010000;
assign label_4[141] = 10'b1000000000;
assign label_4[142] = 10'b1000000000;
assign label_4[143] = 10'b0000010000;
assign label_4[144] = 10'b0010000000;
assign label_4[145] = 10'b0000001000;
assign label_4[146] = 10'b0010000000;
assign label_4[147] = 10'b1000000000;
assign label_4[148] = 10'b1000000000;
assign label_4[149] = 10'b0000000100;
assign label_4[150] = 10'b1000000000;
assign label_4[151] = 10'b0000010000;
assign label_4[152] = 10'b0010000000;
assign label_4[153] = 10'b1000000000;
assign label_4[154] = 10'b0000001000;
assign label_4[155] = 10'b0001000000;
assign label_4[156] = 10'b1000000000;
assign label_4[157] = 10'b0100000000;
assign label_4[158] = 10'b0100000000;
assign label_4[159] = 10'b0000010000;
assign label_4[160] = 10'b0010000000;
assign label_4[161] = 10'b0010000000;
assign label_4[162] = 10'b0000010000;
assign label_4[163] = 10'b0000000100;
assign label_4[164] = 10'b0000001000;
assign label_4[165] = 10'b0010000000;
assign label_4[166] = 10'b0010000000;
assign label_4[167] = 10'b1000000000;
assign label_4[168] = 10'b0000100000;
assign label_4[169] = 10'b0010000000;
assign label_4[170] = 10'b0000000010;
assign label_4[171] = 10'b0000001000;
assign label_4[172] = 10'b0000000100;
assign label_4[173] = 10'b0001000000;
assign label_4[174] = 10'b0000000100;
assign label_4[175] = 10'b0000010000;
assign label_4[176] = 10'b0010000000;
assign label_4[177] = 10'b0010000000;
assign label_4[178] = 10'b1000000000;
assign label_4[179] = 10'b0000000100;
assign label_4[180] = 10'b0010000000;
assign label_4[181] = 10'b0000001000;
assign label_4[182] = 10'b1000000000;
assign label_4[183] = 10'b0010000000;
assign label_4[184] = 10'b0000001000;
assign label_4[185] = 10'b1000000000;
assign label_4[186] = 10'b1000000000;
assign label_4[187] = 10'b0100000000;
assign label_4[188] = 10'b1000000000;
assign label_4[189] = 10'b0010000000;
assign label_4[190] = 10'b0010000000;
assign label_4[191] = 10'b0000001000;
assign label_4[192] = 10'b0000100000;
assign label_4[193] = 10'b0000000100;
assign label_4[194] = 10'b1000000000;
assign label_4[195] = 10'b0000000100;
assign label_4[196] = 10'b0010000000;
assign label_4[197] = 10'b1000000000;
assign label_4[198] = 10'b0000001000;
assign label_4[199] = 10'b0100000000;
assign label_4[200] = 10'b0000100000;
assign label_4[201] = 10'b0000100000;
assign label_4[202] = 10'b0000001000;
assign label_4[203] = 10'b0000000100;
assign label_4[204] = 10'b0100000000;
assign label_4[205] = 10'b0100000000;
assign label_4[206] = 10'b0001000000;
assign label_4[207] = 10'b0000001000;
assign label_4[208] = 10'b0001000000;
assign label_4[209] = 10'b0000010000;
assign label_4[210] = 10'b0000010000;
assign label_4[211] = 10'b0001000000;
assign label_4[212] = 10'b0000000100;
assign label_4[213] = 10'b0000000001;
assign label_4[214] = 10'b0000000100;
assign label_4[215] = 10'b1000000000;
assign label_4[216] = 10'b0100000000;
assign label_4[217] = 10'b0000000100;
assign label_4[218] = 10'b0000010000;
assign label_4[219] = 10'b0000010000;
assign label_4[220] = 10'b0000000100;
assign label_4[221] = 10'b0000000100;
assign label_4[222] = 10'b0010000000;
assign label_4[223] = 10'b0010000000;
assign label_4[224] = 10'b0000100000;
assign label_4[225] = 10'b0000000100;
assign label_4[226] = 10'b0010000000;
assign label_4[227] = 10'b0010000000;
assign label_4[228] = 10'b0000100000;
assign label_4[229] = 10'b0010000000;
assign label_4[230] = 10'b0000000100;
assign label_4[231] = 10'b0000000100;
assign label_4[232] = 10'b0000001000;
assign label_4[233] = 10'b0000001000;
assign label_4[234] = 10'b0100000000;
assign label_4[235] = 10'b0100000000;
assign label_4[236] = 10'b0000001000;
assign label_4[237] = 10'b0000001000;
assign label_4[238] = 10'b0000100000;
assign label_4[239] = 10'b0000001000;
assign label_4[240] = 10'b0001000000;
assign label_4[241] = 10'b0001000000;
assign label_4[242] = 10'b0000000001;
assign label_4[243] = 10'b0000000001;
assign label_4[244] = 10'b0100000000;
assign label_4[245] = 10'b0000000100;
assign label_4[246] = 10'b0100000000;
assign label_4[247] = 10'b0100000000;
assign label_4[248] = 10'b0000000010;
assign label_4[249] = 10'b0000000100;
assign label_4[250] = 10'b0000000100;
assign label_4[251] = 10'b0000001000;
assign label_4[252] = 10'b0000000010;
assign label_4[253] = 10'b0100000000;
assign label_4[254] = 10'b0100000000;
assign label_4[255] = 10'b0100000000;
assign label_4[256] = 10'b0000010000;
assign label_4[257] = 10'b0010000000;
assign label_4[258] = 10'b0000010000;
assign label_4[259] = 10'b1000000000;
assign label_4[260] = 10'b0000010000;
assign label_4[261] = 10'b0000010000;
assign label_4[262] = 10'b1000000000;
assign label_4[263] = 10'b0010000000;
assign label_4[264] = 10'b0000100000;
assign label_4[265] = 10'b0000100000;
assign label_4[266] = 10'b0000100000;
assign label_4[267] = 10'b0000000001;
assign label_4[268] = 10'b0000100000;
assign label_4[269] = 10'b0100000000;
assign label_4[270] = 10'b0000010000;
assign label_4[271] = 10'b1000000000;
assign label_4[272] = 10'b0010000000;
assign label_4[273] = 10'b0000010000;
assign label_4[274] = 10'b0010000000;
assign label_4[275] = 10'b1000000000;
assign label_4[276] = 10'b0000010000;
assign label_4[277] = 10'b1000000000;
assign label_4[278] = 10'b1000000000;
assign label_4[279] = 10'b0000010000;
assign label_4[280] = 10'b0000010000;
assign label_4[281] = 10'b0000010000;
assign label_4[282] = 10'b0000010000;
assign label_4[283] = 10'b0000010000;
assign label_4[284] = 10'b1000000000;
assign label_4[285] = 10'b0010000000;
assign label_4[286] = 10'b0000100000;
assign label_4[287] = 10'b0000010000;
assign label_4[288] = 10'b0000000001;
assign label_4[289] = 10'b0000100000;
assign label_4[290] = 10'b0000010000;
assign label_4[291] = 10'b0010000000;
assign label_4[292] = 10'b0010000000;
assign label_4[293] = 10'b1000000000;
assign label_4[294] = 10'b1000000000;
assign label_4[295] = 10'b1000000000;
assign label_4[296] = 10'b0000010000;
assign label_4[297] = 10'b0000010000;
assign label_4[298] = 10'b1000000000;
assign label_4[299] = 10'b0000010000;
assign label_4[300] = 10'b0100000000;
assign label_4[301] = 10'b0001000000;
assign label_4[302] = 10'b0000010000;
assign label_4[303] = 10'b0001000000;
assign label_4[304] = 10'b0001000000;
assign label_4[305] = 10'b0000000001;
assign label_4[306] = 10'b1000000000;
assign label_4[307] = 10'b0010000000;
assign label_4[308] = 10'b0000001000;
assign label_4[309] = 10'b0000000001;
assign label_4[310] = 10'b0100000000;
assign label_4[311] = 10'b0001000000;
assign label_4[312] = 10'b0000100000;
assign label_4[313] = 10'b0000000001;
assign label_4[314] = 10'b0000000001;
assign label_4[315] = 10'b0100000000;
assign label_4[316] = 10'b0000010000;
assign label_4[317] = 10'b0000100000;
assign label_4[318] = 10'b0001000000;
assign label_4[319] = 10'b0001000000;
assign label_4[320] = 10'b1000000000;
assign label_4[321] = 10'b1000000000;
assign label_4[322] = 10'b0000000001;
assign label_4[323] = 10'b0001000000;
assign label_4[324] = 10'b1000000000;
assign label_4[325] = 10'b1000000000;
assign label_4[326] = 10'b0000000100;
assign label_4[327] = 10'b0000000100;
assign label_4[328] = 10'b0000000001;
assign label_4[329] = 10'b0000100000;
assign label_4[330] = 10'b0000001000;
assign label_4[331] = 10'b0000000100;
assign label_4[332] = 10'b0000000100;
assign label_4[333] = 10'b0000010000;
assign label_4[334] = 10'b1000000000;
assign label_4[335] = 10'b0010000000;
assign label_4[336] = 10'b0000010000;
assign label_4[337] = 10'b1000000000;
assign label_4[338] = 10'b0000001000;
assign label_4[339] = 10'b0000010000;
assign label_4[340] = 10'b0000001000;
assign label_4[341] = 10'b0000001000;
assign label_4[342] = 10'b0000100000;
assign label_4[343] = 10'b0000000001;
assign label_4[344] = 10'b0001000000;
assign label_4[345] = 10'b0000001000;
assign label_4[346] = 10'b0000001000;
assign label_4[347] = 10'b0000100000;
assign label_4[348] = 10'b1000000000;
assign label_4[349] = 10'b0000000001;
assign label_4[350] = 10'b0000001000;
assign label_4[351] = 10'b0100000000;
assign label_4[352] = 10'b0000100000;
assign label_4[353] = 10'b0000000001;
assign label_4[354] = 10'b0000100000;
assign label_4[355] = 10'b0000100000;
assign label_4[356] = 10'b0000100000;
assign label_4[357] = 10'b0100000000;
assign label_4[358] = 10'b0000001000;
assign label_4[359] = 10'b0100000000;
assign label_4[360] = 10'b0000000100;
assign label_4[361] = 10'b0000000100;
assign label_4[362] = 10'b0000000100;
assign label_4[363] = 10'b0000000100;
assign label_4[364] = 10'b0000000100;
assign label_4[365] = 10'b0000000100;
assign label_4[366] = 10'b0001000000;
assign label_4[367] = 10'b0000000001;
assign label_4[368] = 10'b0000010000;
assign label_4[369] = 10'b0000010000;
assign label_4[370] = 10'b0000000100;
assign label_4[371] = 10'b0000000001;
assign label_4[372] = 10'b0000000100;
assign label_4[373] = 10'b0000000100;
assign label_4[374] = 10'b0000000001;
assign label_4[375] = 10'b0000001000;
assign label_4[376] = 10'b1000000000;
assign label_4[377] = 10'b1000000000;
assign label_4[378] = 10'b0000001000;
assign label_4[379] = 10'b1000000000;
assign label_4[380] = 10'b1000000000;
assign label_4[381] = 10'b0000000100;
assign label_4[382] = 10'b0100000000;
assign label_4[383] = 10'b0000000100;
assign label_4[384] = 10'b1000000000;
assign label_4[385] = 10'b0100000000;
assign label_4[386] = 10'b0000100000;
assign label_4[387] = 10'b1000000000;
assign label_4[388] = 10'b0000000001;
assign label_4[389] = 10'b0000000001;
assign label_4[390] = 10'b0000000001;
assign label_4[391] = 10'b0000000001;
assign label_4[392] = 10'b0000100000;
assign label_4[393] = 10'b0000100000;
assign label_4[394] = 10'b0000100000;
assign label_4[395] = 10'b0000100000;
assign label_4[396] = 10'b0000100000;
assign label_4[397] = 10'b0100000000;
assign label_4[398] = 10'b0100000000;
assign label_4[399] = 10'b0100000000;
assign label_4[400] = 10'b0000010000;
assign label_4[401] = 10'b0100000000;
assign label_4[402] = 10'b0100000000;
assign label_4[403] = 10'b0100000000;
assign label_4[404] = 10'b0000010000;
assign label_4[405] = 10'b0000010000;
assign label_4[406] = 10'b0010000000;
assign label_4[407] = 10'b0010000000;
assign label_4[408] = 10'b0100000000;
assign label_4[409] = 10'b0100000000;
assign label_4[410] = 10'b0100000000;
assign label_4[411] = 10'b0100000000;
assign label_4[412] = 10'b0010000000;
assign label_4[413] = 10'b1000000000;
assign label_4[414] = 10'b0100000000;
assign label_4[415] = 10'b0000010000;
assign label_4[416] = 10'b0000100000;
assign label_4[417] = 10'b0000100000;
assign label_4[418] = 10'b0000100000;
assign label_4[419] = 10'b0100000000;
assign label_4[420] = 10'b0000100000;
assign label_4[421] = 10'b0000100000;
assign label_4[422] = 10'b0000100000;
assign label_4[423] = 10'b0100000000;
assign label_4[424] = 10'b0000000001;
assign label_4[425] = 10'b0000100000;
assign label_4[426] = 10'b0000000001;
assign label_4[427] = 10'b0000010000;
assign label_4[428] = 10'b0000100000;
assign label_4[429] = 10'b0000100000;
assign label_4[430] = 10'b0100000000;
assign label_4[431] = 10'b0100000000;
assign label_4[432] = 10'b0010000000;
assign label_4[433] = 10'b0010000000;
assign label_4[434] = 10'b0010000000;
assign label_4[435] = 10'b0010000000;
assign label_4[436] = 10'b1000000000;
assign label_4[437] = 10'b1000000000;
assign label_4[438] = 10'b0010000000;
assign label_4[439] = 10'b1000000000;
assign label_4[440] = 10'b0010000000;
assign label_4[441] = 10'b0010000000;
assign label_4[442] = 10'b0010000000;
assign label_4[443] = 10'b0010000000;
assign label_4[444] = 10'b0010000000;
assign label_4[445] = 10'b0010000000;
assign label_4[446] = 10'b0010000000;
assign label_4[447] = 10'b0010000000;
assign label_4[448] = 10'b0001000000;
assign label_4[449] = 10'b0000100000;
assign label_4[450] = 10'b0000000001;
assign label_4[451] = 10'b0000100000;
assign label_4[452] = 10'b0100000000;
assign label_4[453] = 10'b0000010000;
assign label_4[454] = 10'b0000010000;
assign label_4[455] = 10'b0000001000;
assign label_4[456] = 10'b0001000000;
assign label_4[457] = 10'b0001000000;
assign label_4[458] = 10'b0001000000;
assign label_4[459] = 10'b0001000000;
assign label_4[460] = 10'b0001000000;
assign label_4[461] = 10'b0001000000;
assign label_4[462] = 10'b0001000000;
assign label_4[463] = 10'b0001000000;
assign label_4[464] = 10'b0000100000;
assign label_4[465] = 10'b0000010000;
assign label_4[466] = 10'b0100000000;
assign label_4[467] = 10'b0000010000;
assign label_4[468] = 10'b0000010000;
assign label_4[469] = 10'b0001000000;
assign label_4[470] = 10'b0000010000;
assign label_4[471] = 10'b0010000000;
assign label_4[472] = 10'b0100000000;
assign label_4[473] = 10'b0010000000;
assign label_4[474] = 10'b1000000000;
assign label_4[475] = 10'b1000000000;
assign label_4[476] = 10'b0100000000;
assign label_4[477] = 10'b0000100000;
assign label_4[478] = 10'b0100000000;
assign label_4[479] = 10'b0000100000;
assign label_4[480] = 10'b0000000100;
assign label_4[481] = 10'b0000010000;
assign label_4[482] = 10'b0100000000;
assign label_4[483] = 10'b0000000100;
assign label_4[484] = 10'b0000100000;
assign label_4[485] = 10'b0000100000;
assign label_4[486] = 10'b0100000000;
assign label_4[487] = 10'b0100000000;
assign label_4[488] = 10'b0000000001;
assign label_4[489] = 10'b0000100000;
assign label_4[490] = 10'b0001000000;
assign label_4[491] = 10'b0000001000;
assign label_4[492] = 10'b0001000000;
assign label_4[493] = 10'b0000010000;
assign label_4[494] = 10'b0100000000;
assign label_4[495] = 10'b0100000000;
assign label_4[496] = 10'b0000000001;
assign label_4[497] = 10'b0000100000;
assign label_4[498] = 10'b0000100000;
assign label_4[499] = 10'b0000100000;
assign label_4[500] = 10'b0000000001;
assign label_4[501] = 10'b0000000001;
assign label_4[502] = 10'b0001000000;
assign label_4[503] = 10'b0000000001;
assign label_4[504] = 10'b0000100000;
assign label_4[505] = 10'b0000000001;
assign label_4[506] = 10'b0000000001;
assign label_4[507] = 10'b0100000000;
assign label_4[508] = 10'b0000010000;
assign label_4[509] = 10'b0000000001;
assign label_4[510] = 10'b0100000000;
assign label_4[511] = 10'b0000000001;
assign label_4[512] = 10'b0000000100;
assign label_4[513] = 10'b0000100000;
assign label_4[514] = 10'b0000001000;
assign label_4[515] = 10'b0000000100;
assign label_4[516] = 10'b0000000001;
assign label_4[517] = 10'b0000000001;
assign label_4[518] = 10'b0000000100;
assign label_4[519] = 10'b0000100000;
assign label_4[520] = 10'b0000010000;
assign label_4[521] = 10'b0000000100;
assign label_4[522] = 10'b0100000000;
assign label_4[523] = 10'b0000001000;
assign label_4[524] = 10'b0000000100;
assign label_4[525] = 10'b0000001000;
assign label_4[526] = 10'b0000000100;
assign label_4[527] = 10'b0100000000;
assign label_4[528] = 10'b0000000010;
assign label_4[529] = 10'b0000010000;
assign label_4[530] = 10'b0000001000;
assign label_4[531] = 10'b0000010000;
assign label_4[532] = 10'b0000001000;
assign label_4[533] = 10'b0000100000;
assign label_4[534] = 10'b0000001000;
assign label_4[535] = 10'b0100000000;
assign label_4[536] = 10'b0000001000;
assign label_4[537] = 10'b0000000100;
assign label_4[538] = 10'b0000000100;
assign label_4[539] = 10'b0000001000;
assign label_4[540] = 10'b0000010000;
assign label_4[541] = 10'b0100000000;
assign label_4[542] = 10'b0000000100;
assign label_4[543] = 10'b0000100000;
assign label_4[544] = 10'b0000001000;
assign label_4[545] = 10'b0001000000;
assign label_4[546] = 10'b0000100000;
assign label_4[547] = 10'b0001000000;
assign label_4[548] = 10'b0100000000;
assign label_4[549] = 10'b0100000000;
assign label_4[550] = 10'b0000000001;
assign label_4[551] = 10'b0000010000;
assign label_4[552] = 10'b0000000001;
assign label_4[553] = 10'b0100000000;
assign label_4[554] = 10'b0000000001;
assign label_4[555] = 10'b0000000001;
assign label_4[556] = 10'b0000000001;
assign label_4[557] = 10'b0100000000;
assign label_4[558] = 10'b0100000000;
assign label_4[559] = 10'b0100000000;
assign label_4[560] = 10'b0000100000;
assign label_4[561] = 10'b0100000000;
assign label_4[562] = 10'b0100000000;
assign label_4[563] = 10'b0000000001;
assign label_4[564] = 10'b0000000001;
assign label_4[565] = 10'b0000010000;
assign label_4[566] = 10'b0100000000;
assign label_4[567] = 10'b0001000000;
assign label_4[568] = 10'b0000001000;
assign label_4[569] = 10'b0100000000;
assign label_4[570] = 10'b0100000000;
assign label_4[571] = 10'b0100000000;
assign label_4[572] = 10'b0000001000;
assign label_4[573] = 10'b0000001000;
assign label_4[574] = 10'b0000000100;
assign label_4[575] = 10'b0000000100;
assign label_4[576] = 10'b0000100000;
assign label_4[577] = 10'b0000000100;
assign label_4[578] = 10'b0000000001;
assign label_4[579] = 10'b0000100000;
assign label_4[580] = 10'b0001000000;
assign label_4[581] = 10'b0000000001;
assign label_4[582] = 10'b0000000001;
assign label_4[583] = 10'b0000100000;
assign label_4[584] = 10'b0000000001;
assign label_4[585] = 10'b0000000001;
assign label_4[586] = 10'b0000000001;
assign label_4[587] = 10'b0000100000;
assign label_4[588] = 10'b0000100000;
assign label_4[589] = 10'b0000010000;
assign label_4[590] = 10'b0000000100;
assign label_4[591] = 10'b0000000100;
assign label_4[592] = 10'b0000100000;
assign label_4[593] = 10'b0000100000;
assign label_4[594] = 10'b0000010000;
assign label_4[595] = 10'b0100000000;
assign label_4[596] = 10'b0100000000;
assign label_4[597] = 10'b0100000000;
assign label_4[598] = 10'b0100000000;
assign label_4[599] = 10'b0000100000;
assign label_4[600] = 10'b0000100000;
assign label_4[601] = 10'b0000100000;
assign label_4[602] = 10'b0000100000;
assign label_4[603] = 10'b0000100000;
assign label_4[604] = 10'b0000100000;
assign label_4[605] = 10'b0001000000;
assign label_4[606] = 10'b0000100000;
assign label_4[607] = 10'b0001000000;
assign label_4[608] = 10'b0000001000;
assign label_4[609] = 10'b0000100000;
assign label_4[610] = 10'b0000100000;
assign label_4[611] = 10'b0100000000;
assign label_4[612] = 10'b0100000000;
assign label_4[613] = 10'b0100000000;
assign label_4[614] = 10'b0000001000;
assign label_4[615] = 10'b0100000000;
assign label_4[616] = 10'b0000010000;
assign label_4[617] = 10'b0000000100;
assign label_4[618] = 10'b0000010000;
assign label_4[619] = 10'b0100000000;
assign label_4[620] = 10'b0100000000;
assign label_4[621] = 10'b0100000000;
assign label_4[622] = 10'b0000000100;
assign label_4[623] = 10'b0100000000;
assign label_4[624] = 10'b0000100000;
assign label_4[625] = 10'b0000001000;
assign label_4[626] = 10'b0100000000;
assign label_4[627] = 10'b0000001000;
assign label_4[628] = 10'b0100000000;
assign label_4[629] = 10'b0100000000;
assign label_4[630] = 10'b0100000000;
assign label_4[631] = 10'b0000001000;
assign label_4[632] = 10'b0100000000;
assign label_4[633] = 10'b0000000001;
assign label_4[634] = 10'b0000001000;
assign label_4[635] = 10'b0000000001;
assign label_4[636] = 10'b0100000000;
assign label_4[637] = 10'b0100000000;
assign label_4[638] = 10'b0100000000;
assign label_4[639] = 10'b0000001000;
assign label_4[640] = 10'b0000100000;
assign label_4[641] = 10'b0000001000;
assign label_4[642] = 10'b0000001000;
assign label_4[643] = 10'b0000000001;
assign label_4[644] = 10'b0000100000;
assign label_4[645] = 10'b0000001000;
assign label_4[646] = 10'b0000100000;
assign label_4[647] = 10'b0100000000;
assign label_4[648] = 10'b0001000000;
assign label_4[649] = 10'b0001000000;
assign label_4[650] = 10'b0001000000;
assign label_4[651] = 10'b0000100000;
assign label_4[652] = 10'b0000000100;
assign label_4[653] = 10'b0000001000;
assign label_4[654] = 10'b0100000000;
assign label_4[655] = 10'b1000000000;
assign label_4[656] = 10'b0000010000;
assign label_4[657] = 10'b1000000000;
assign label_4[658] = 10'b0000010000;
assign label_4[659] = 10'b0000010000;
assign label_4[660] = 10'b0000000100;
assign label_4[661] = 10'b0000100000;
assign label_4[662] = 10'b0000001000;
assign label_4[663] = 10'b0000001000;
assign label_4[664] = 10'b0000000100;
assign label_4[665] = 10'b0000000100;
assign label_4[666] = 10'b0000010000;
assign label_4[667] = 10'b0001000000;
assign label_4[668] = 10'b0001000000;
assign label_4[669] = 10'b0100000000;
assign label_4[670] = 10'b0100000000;
assign label_4[671] = 10'b0100000000;
assign label_4[672] = 10'b0000000001;
assign label_4[673] = 10'b0000100000;
assign label_4[674] = 10'b0000000001;
assign label_4[675] = 10'b0000000001;
assign label_4[676] = 10'b0100000000;
assign label_4[677] = 10'b0000000001;
assign label_4[678] = 10'b1000000000;
assign label_4[679] = 10'b0000000001;
assign label_4[680] = 10'b0000100000;
assign label_4[681] = 10'b0000001000;
assign label_4[682] = 10'b0000000001;
assign label_4[683] = 10'b0000100000;
assign label_4[684] = 10'b0000001000;
assign label_4[685] = 10'b0000100000;
assign label_4[686] = 10'b0000001000;
assign label_4[687] = 10'b0000001000;
assign label_4[688] = 10'b0000001000;
assign label_4[689] = 10'b0000000001;
assign label_4[690] = 10'b0000000001;
assign label_4[691] = 10'b0000000001;
assign label_4[692] = 10'b0001000000;
assign label_4[693] = 10'b0000000001;
assign label_4[694] = 10'b0100000000;
assign label_4[695] = 10'b0000001000;
assign label_4[696] = 10'b0000010000;
assign label_4[697] = 10'b1000000000;
assign label_4[698] = 10'b0100000000;
assign label_4[699] = 10'b0000001000;
assign label_4[700] = 10'b0000000100;
assign label_4[701] = 10'b0000000100;
assign label_4[702] = 10'b0000000100;
assign label_4[703] = 10'b0000000001;
assign label_4[704] = 10'b0000000100;
assign label_4[705] = 10'b0100000000;
assign label_4[706] = 10'b0000000001;
assign label_4[707] = 10'b0000000001;
assign label_4[708] = 10'b0000000001;
assign label_4[709] = 10'b0000000001;
assign label_4[710] = 10'b0000000001;
assign label_4[711] = 10'b0000000001;
assign label_4[712] = 10'b0000000001;
assign label_4[713] = 10'b0000000001;
assign label_4[714] = 10'b0000000001;
assign label_4[715] = 10'b0000000001;
assign label_4[716] = 10'b0000001000;
assign label_4[717] = 10'b0000000001;
assign label_4[718] = 10'b0100000000;
assign label_4[719] = 10'b0100000000;
assign label_4[720] = 10'b0000000001;
assign label_4[721] = 10'b0000000001;
assign label_4[722] = 10'b0000000001;
assign label_4[723] = 10'b0000000001;
assign label_4[724] = 10'b0000010000;
assign label_4[725] = 10'b0000010000;
assign label_4[726] = 10'b1000000000;
assign label_4[727] = 10'b1000000000;
assign label_4[728] = 10'b0000000001;
assign label_4[729] = 10'b0000000001;
assign label_4[730] = 10'b0000000001;
assign label_4[731] = 10'b0000000001;
assign label_4[732] = 10'b0000000001;
assign label_4[733] = 10'b0000000001;
assign label_4[734] = 10'b0000000001;
assign label_4[735] = 10'b0000000001;
assign label_4[736] = 10'b0100000000;
assign label_4[737] = 10'b0100000000;
assign label_4[738] = 10'b0000001000;
assign label_4[739] = 10'b0000001000;
assign label_4[740] = 10'b0000001000;
assign label_4[741] = 10'b0000001000;
assign label_4[742] = 10'b0000001000;
assign label_4[743] = 10'b0000001000;
assign label_4[744] = 10'b0000000001;
assign label_4[745] = 10'b0000000001;
assign label_4[746] = 10'b0000000001;
assign label_4[747] = 10'b0000000001;
assign label_4[748] = 10'b0000010000;
assign label_4[749] = 10'b0000010000;
assign label_4[750] = 10'b0100000000;
assign label_4[751] = 10'b0100000000;
assign label_4[752] = 10'b0000000100;
assign label_4[753] = 10'b0000000001;
assign label_4[754] = 10'b0000001000;
assign label_4[755] = 10'b0000001000;
assign label_4[756] = 10'b0000000100;
assign label_4[757] = 10'b0000000001;
assign label_4[758] = 10'b1000000000;
assign label_4[759] = 10'b1000000000;
assign label_4[760] = 10'b0000000001;
assign label_4[761] = 10'b0100000000;
assign label_4[762] = 10'b0000000001;
assign label_4[763] = 10'b0000010000;
assign label_4[764] = 10'b0000000001;
assign label_4[765] = 10'b0100000000;
assign label_4[766] = 10'b0000001000;
assign label_4[767] = 10'b0000000001;
assign label_4[768] = 10'b0000000010;
assign label_4[769] = 10'b0000000010;
assign label_4[770] = 10'b0001000000;
assign label_4[771] = 10'b0000000001;
assign label_4[772] = 10'b0010000000;
assign label_4[773] = 10'b0000000010;
assign label_4[774] = 10'b0000000100;
assign label_4[775] = 10'b0000100000;
assign label_4[776] = 10'b0000010000;
assign label_4[777] = 10'b0000000100;
assign label_4[778] = 10'b0000001000;
assign label_4[779] = 10'b0000100000;
assign label_4[780] = 10'b0100000000;
assign label_4[781] = 10'b0000000100;
assign label_4[782] = 10'b0000001000;
assign label_4[783] = 10'b0000000100;
assign label_4[784] = 10'b0000000100;
assign label_4[785] = 10'b0000001000;
assign label_4[786] = 10'b0000001000;
assign label_4[787] = 10'b0001000000;
assign label_4[788] = 10'b0000000010;
assign label_4[789] = 10'b0100000000;
assign label_4[790] = 10'b0000001000;
assign label_4[791] = 10'b0000001000;
assign label_4[792] = 10'b0100000000;
assign label_4[793] = 10'b0100000000;
assign label_4[794] = 10'b0000010000;
assign label_4[795] = 10'b0100000000;
assign label_4[796] = 10'b0000000010;
assign label_4[797] = 10'b0000100000;
assign label_4[798] = 10'b1000000000;
assign label_4[799] = 10'b0000001000;
assign label_4[800] = 10'b0000000100;
assign label_4[801] = 10'b0000000100;
assign label_4[802] = 10'b0001000000;
assign label_4[803] = 10'b0001000000;
assign label_4[804] = 10'b0010000000;
assign label_4[805] = 10'b0000001000;
assign label_4[806] = 10'b0000000100;
assign label_4[807] = 10'b0000001000;
assign label_4[808] = 10'b0001000000;
assign label_4[809] = 10'b0100000000;
assign label_4[810] = 10'b0100000000;
assign label_4[811] = 10'b0000000001;
assign label_4[812] = 10'b0000001000;
assign label_4[813] = 10'b0000001000;
assign label_4[814] = 10'b0000000001;
assign label_4[815] = 10'b0000000100;
assign label_4[816] = 10'b0000010000;
assign label_4[817] = 10'b0001000000;
assign label_4[818] = 10'b0000010000;
assign label_4[819] = 10'b0000010000;
assign label_4[820] = 10'b0001000000;
assign label_4[821] = 10'b0000010000;
assign label_4[822] = 10'b0001000000;
assign label_4[823] = 10'b0000000100;
assign label_4[824] = 10'b0000000001;
assign label_4[825] = 10'b0000100000;
assign label_4[826] = 10'b0000000100;
assign label_4[827] = 10'b0100000000;
assign label_4[828] = 10'b0000000001;
assign label_4[829] = 10'b0001000000;
assign label_4[830] = 10'b0000100000;
assign label_4[831] = 10'b0001000000;
assign label_4[832] = 10'b0000000100;
assign label_4[833] = 10'b0000000100;
assign label_4[834] = 10'b0000000010;
assign label_4[835] = 10'b0100000000;
assign label_4[836] = 10'b0100000000;
assign label_4[837] = 10'b0100000000;
assign label_4[838] = 10'b0000100000;
assign label_4[839] = 10'b0000000100;
assign label_4[840] = 10'b0001000000;
assign label_4[841] = 10'b0000000100;
assign label_4[842] = 10'b0000000010;
assign label_4[843] = 10'b0000000100;
assign label_4[844] = 10'b0000000100;
assign label_4[845] = 10'b0100000000;
assign label_4[846] = 10'b0000000100;
assign label_4[847] = 10'b0100000000;
assign label_4[848] = 10'b0000000100;
assign label_4[849] = 10'b0000000100;
assign label_4[850] = 10'b0010000000;
assign label_4[851] = 10'b0100000000;
assign label_4[852] = 10'b1000000000;
assign label_4[853] = 10'b0001000000;
assign label_4[854] = 10'b0100000000;
assign label_4[855] = 10'b0100000000;
assign label_4[856] = 10'b0100000000;
assign label_4[857] = 10'b0000000100;
assign label_4[858] = 10'b0001000000;
assign label_4[859] = 10'b0000000100;
assign label_4[860] = 10'b0000000100;
assign label_4[861] = 10'b0000000100;
assign label_4[862] = 10'b0100000000;
assign label_4[863] = 10'b0000000100;
assign label_4[864] = 10'b0001000000;
assign label_4[865] = 10'b0000010000;
assign label_4[866] = 10'b0001000000;
assign label_4[867] = 10'b0000000001;
assign label_4[868] = 10'b0000010000;
assign label_4[869] = 10'b0010000000;
assign label_4[870] = 10'b0000000001;
assign label_4[871] = 10'b0100000000;
assign label_4[872] = 10'b0000100000;
assign label_4[873] = 10'b0000000100;
assign label_4[874] = 10'b0000000001;
assign label_4[875] = 10'b0000000001;
assign label_4[876] = 10'b0100000000;
assign label_4[877] = 10'b0100000000;
assign label_4[878] = 10'b0000000100;
assign label_4[879] = 10'b0000010000;
assign label_4[880] = 10'b0000100000;
assign label_4[881] = 10'b0100000000;
assign label_4[882] = 10'b0000010000;
assign label_4[883] = 10'b0000010000;
assign label_4[884] = 10'b0100000000;
assign label_4[885] = 10'b0100000000;
assign label_4[886] = 10'b0000010000;
assign label_4[887] = 10'b0100000000;
assign label_4[888] = 10'b1000000000;
assign label_4[889] = 10'b1000000000;
assign label_4[890] = 10'b1000000000;
assign label_4[891] = 10'b1000000000;
assign label_4[892] = 10'b0100000000;
assign label_4[893] = 10'b0100000000;
assign label_4[894] = 10'b0000010000;
assign label_4[895] = 10'b0000000001;
assign label_4[896] = 10'b0000000100;
assign label_4[897] = 10'b0000000100;
assign label_4[898] = 10'b0100000000;
assign label_4[899] = 10'b0000100000;
assign label_4[900] = 10'b0000000100;
assign label_4[901] = 10'b0000000100;
assign label_4[902] = 10'b1000000000;
assign label_4[903] = 10'b0000000100;
assign label_4[904] = 10'b0010000000;
assign label_4[905] = 10'b0100000000;
assign label_4[906] = 10'b0100000000;
assign label_4[907] = 10'b0100000000;
assign label_4[908] = 10'b0000000001;
assign label_4[909] = 10'b0100000000;
assign label_4[910] = 10'b0000000100;
assign label_4[911] = 10'b0000000100;
assign label_4[912] = 10'b0000000010;
assign label_4[913] = 10'b0000001000;
assign label_4[914] = 10'b0100000000;
assign label_4[915] = 10'b0000001000;
assign label_4[916] = 10'b0000001000;
assign label_4[917] = 10'b0100000000;
assign label_4[918] = 10'b0000000001;
assign label_4[919] = 10'b0100000000;
assign label_4[920] = 10'b0000100000;
assign label_4[921] = 10'b0000001000;
assign label_4[922] = 10'b0000001000;
assign label_4[923] = 10'b0000001000;
assign label_4[924] = 10'b0000100000;
assign label_4[925] = 10'b0000100000;
assign label_4[926] = 10'b0100000000;
assign label_4[927] = 10'b0100000000;
assign label_4[928] = 10'b0000000100;
assign label_4[929] = 10'b0000000100;
assign label_4[930] = 10'b0000000100;
assign label_4[931] = 10'b0000000100;
assign label_4[932] = 10'b0000000100;
assign label_4[933] = 10'b0100000000;
assign label_4[934] = 10'b0000000100;
assign label_4[935] = 10'b0000000001;
assign label_4[936] = 10'b0000000001;
assign label_4[937] = 10'b0000000100;
assign label_4[938] = 10'b0000000001;
assign label_4[939] = 10'b0000000100;
assign label_4[940] = 10'b0000000100;
assign label_4[941] = 10'b0000000100;
assign label_4[942] = 10'b0000000001;
assign label_4[943] = 10'b1000000000;
assign label_4[944] = 10'b0000000010;
assign label_4[945] = 10'b0000000100;
assign label_4[946] = 10'b0000001000;
assign label_4[947] = 10'b0000001000;
assign label_4[948] = 10'b0000001000;
assign label_4[949] = 10'b0100000000;
assign label_4[950] = 10'b0100000000;
assign label_4[951] = 10'b0100000000;
assign label_4[952] = 10'b0000000100;
assign label_4[953] = 10'b0000000100;
assign label_4[954] = 10'b0000001000;
assign label_4[955] = 10'b0000001000;
assign label_4[956] = 10'b0000001000;
assign label_4[957] = 10'b0000100000;
assign label_4[958] = 10'b0000000100;
assign label_4[959] = 10'b0000000100;
assign label_4[960] = 10'b0000000001;
assign label_4[961] = 10'b0000010000;
assign label_4[962] = 10'b0100000000;
assign label_4[963] = 10'b1000000000;
assign label_4[964] = 10'b0000000100;
assign label_4[965] = 10'b0000000100;
assign label_4[966] = 10'b0000000001;
assign label_4[967] = 10'b1000000000;
assign label_4[968] = 10'b0000000100;
assign label_4[969] = 10'b0000000001;
assign label_4[970] = 10'b0000000100;
assign label_4[971] = 10'b0000000100;
assign label_4[972] = 10'b0000000001;
assign label_4[973] = 10'b0000000001;
assign label_4[974] = 10'b0000100000;
assign label_4[975] = 10'b0000100000;
assign label_4[976] = 10'b0000001000;
assign label_4[977] = 10'b0000001000;
assign label_4[978] = 10'b0000000001;
assign label_4[979] = 10'b0000001000;
assign label_4[980] = 10'b0000000001;
assign label_4[981] = 10'b0000001000;
assign label_4[982] = 10'b0000000001;
assign label_4[983] = 10'b0000000001;
assign label_4[984] = 10'b0000001000;
assign label_4[985] = 10'b0000000100;
assign label_4[986] = 10'b0100000000;
assign label_4[987] = 10'b0000001000;
assign label_4[988] = 10'b0100000000;
assign label_4[989] = 10'b0000000001;
assign label_4[990] = 10'b0000000100;
assign label_4[991] = 10'b0000000001;
assign label_4[992] = 10'b0100000000;
assign label_4[993] = 10'b1000000000;
assign label_4[994] = 10'b0000100000;
assign label_4[995] = 10'b0000000100;
assign label_4[996] = 10'b0000000100;
assign label_4[997] = 10'b0000000001;
assign label_4[998] = 10'b0001000000;
assign label_4[999] = 10'b0000000100;
assign label_4[1000] = 10'b0000001000;
assign label_4[1001] = 10'b0100000000;
assign label_4[1002] = 10'b0000100000;
assign label_4[1003] = 10'b0100000000;
assign label_4[1004] = 10'b0000010000;
assign label_4[1005] = 10'b0000000001;
assign label_4[1006] = 10'b0000001000;
assign label_4[1007] = 10'b0000000001;
assign label_4[1008] = 10'b0000000100;
assign label_4[1009] = 10'b0000000100;
assign label_4[1010] = 10'b0001000000;
assign label_4[1011] = 10'b0100000000;
assign label_4[1012] = 10'b0000000100;
assign label_4[1013] = 10'b0100000000;
assign label_4[1014] = 10'b0100000000;
assign label_4[1015] = 10'b0000001000;
assign label_4[1016] = 10'b0000000001;
assign label_4[1017] = 10'b0000000100;
assign label_4[1018] = 10'b0000000001;
assign label_4[1019] = 10'b0100000000;
assign label_4[1020] = 10'b0000000100;
assign label_4[1021] = 10'b0000000100;
assign label_4[1022] = 10'b0000001000;
assign label_4[1023] = 10'b0000001000;
assign label_5[0] = 10'b0000100000;
assign label_5[1] = 10'b0000000001;
assign label_5[2] = 10'b0000000001;
assign label_5[3] = 10'b0010000000;
assign label_5[4] = 10'b0010000000;
assign label_5[5] = 10'b0000010000;
assign label_5[6] = 10'b0010000000;
assign label_5[7] = 10'b0000100000;
assign label_5[8] = 10'b0000100000;
assign label_5[9] = 10'b0000100000;
assign label_5[10] = 10'b0000100000;
assign label_5[11] = 10'b0000000001;
assign label_5[12] = 10'b0000000001;
assign label_5[13] = 10'b0000100000;
assign label_5[14] = 10'b0000000001;
assign label_5[15] = 10'b0000000001;
assign label_5[16] = 10'b0000000001;
assign label_5[17] = 10'b0000000001;
assign label_5[18] = 10'b0000000100;
assign label_5[19] = 10'b0000000001;
assign label_5[20] = 10'b0000100000;
assign label_5[21] = 10'b0000100000;
assign label_5[22] = 10'b0001000000;
assign label_5[23] = 10'b0001000000;
assign label_5[24] = 10'b0000001000;
assign label_5[25] = 10'b0000100000;
assign label_5[26] = 10'b0000100000;
assign label_5[27] = 10'b0000000001;
assign label_5[28] = 10'b0000000001;
assign label_5[29] = 10'b0000001000;
assign label_5[30] = 10'b0000000001;
assign label_5[31] = 10'b0000000001;
assign label_5[32] = 10'b0010000000;
assign label_5[33] = 10'b1000000000;
assign label_5[34] = 10'b0010000000;
assign label_5[35] = 10'b0000000100;
assign label_5[36] = 10'b0000000001;
assign label_5[37] = 10'b0001000000;
assign label_5[38] = 10'b1000000000;
assign label_5[39] = 10'b0000000100;
assign label_5[40] = 10'b0010000000;
assign label_5[41] = 10'b0000100000;
assign label_5[42] = 10'b0000001000;
assign label_5[43] = 10'b0000100000;
assign label_5[44] = 10'b0010000000;
assign label_5[45] = 10'b0010000000;
assign label_5[46] = 10'b0000100000;
assign label_5[47] = 10'b0000001000;
assign label_5[48] = 10'b0000100000;
assign label_5[49] = 10'b0001000000;
assign label_5[50] = 10'b0010000000;
assign label_5[51] = 10'b1000000000;
assign label_5[52] = 10'b0000010000;
assign label_5[53] = 10'b0000010000;
assign label_5[54] = 10'b1000000000;
assign label_5[55] = 10'b0000000001;
assign label_5[56] = 10'b0001000000;
assign label_5[57] = 10'b0010000000;
assign label_5[58] = 10'b1000000000;
assign label_5[59] = 10'b0000010000;
assign label_5[60] = 10'b0000000001;
assign label_5[61] = 10'b0000010000;
assign label_5[62] = 10'b0000000001;
assign label_5[63] = 10'b0000000001;
assign label_5[64] = 10'b0000100000;
assign label_5[65] = 10'b0000100000;
assign label_5[66] = 10'b0000100000;
assign label_5[67] = 10'b0001000000;
assign label_5[68] = 10'b0000010000;
assign label_5[69] = 10'b0000000001;
assign label_5[70] = 10'b0000001000;
assign label_5[71] = 10'b0001000000;
assign label_5[72] = 10'b0001000000;
assign label_5[73] = 10'b0001000000;
assign label_5[74] = 10'b0001000000;
assign label_5[75] = 10'b0001000000;
assign label_5[76] = 10'b0000000100;
assign label_5[77] = 10'b0000000100;
assign label_5[78] = 10'b0000000100;
assign label_5[79] = 10'b0000000100;
assign label_5[80] = 10'b0000010000;
assign label_5[81] = 10'b0000000100;
assign label_5[82] = 10'b1000000000;
assign label_5[83] = 10'b0010000000;
assign label_5[84] = 10'b0000010000;
assign label_5[85] = 10'b0000010000;
assign label_5[86] = 10'b0000100000;
assign label_5[87] = 10'b1000000000;
assign label_5[88] = 10'b0000000100;
assign label_5[89] = 10'b0001000000;
assign label_5[90] = 10'b0000010000;
assign label_5[91] = 10'b0001000000;
assign label_5[92] = 10'b0000000100;
assign label_5[93] = 10'b0100000000;
assign label_5[94] = 10'b0000000001;
assign label_5[95] = 10'b0000100000;
assign label_5[96] = 10'b0000100000;
assign label_5[97] = 10'b0100000000;
assign label_5[98] = 10'b0000100000;
assign label_5[99] = 10'b0000100000;
assign label_5[100] = 10'b0000000100;
assign label_5[101] = 10'b0000000100;
assign label_5[102] = 10'b0000000001;
assign label_5[103] = 10'b0000000001;
assign label_5[104] = 10'b0000000001;
assign label_5[105] = 10'b0000000001;
assign label_5[106] = 10'b0000000001;
assign label_5[107] = 10'b0000000001;
assign label_5[108] = 10'b0000000100;
assign label_5[109] = 10'b0000000100;
assign label_5[110] = 10'b0000100000;
assign label_5[111] = 10'b0000100000;
assign label_5[112] = 10'b0000000100;
assign label_5[113] = 10'b0000000100;
assign label_5[114] = 10'b0000000001;
assign label_5[115] = 10'b0000000001;
assign label_5[116] = 10'b0100000000;
assign label_5[117] = 10'b0100000000;
assign label_5[118] = 10'b0000010000;
assign label_5[119] = 10'b0000000100;
assign label_5[120] = 10'b0000100000;
assign label_5[121] = 10'b0000100000;
assign label_5[122] = 10'b0000000001;
assign label_5[123] = 10'b0000000001;
assign label_5[124] = 10'b1000000000;
assign label_5[125] = 10'b1000000000;
assign label_5[126] = 10'b0000000001;
assign label_5[127] = 10'b0000000001;
assign label_5[128] = 10'b0000001000;
assign label_5[129] = 10'b0000100000;
assign label_5[130] = 10'b0000001000;
assign label_5[131] = 10'b0000100000;
assign label_5[132] = 10'b0000100000;
assign label_5[133] = 10'b0000000001;
assign label_5[134] = 10'b0000001000;
assign label_5[135] = 10'b0000000001;
assign label_5[136] = 10'b0000100000;
assign label_5[137] = 10'b0000001000;
assign label_5[138] = 10'b0000100000;
assign label_5[139] = 10'b0000000001;
assign label_5[140] = 10'b0000100000;
assign label_5[141] = 10'b0000100000;
assign label_5[142] = 10'b0000000100;
assign label_5[143] = 10'b0000000100;
assign label_5[144] = 10'b0000000100;
assign label_5[145] = 10'b0000001000;
assign label_5[146] = 10'b0000100000;
assign label_5[147] = 10'b0000100000;
assign label_5[148] = 10'b0000000100;
assign label_5[149] = 10'b0000000100;
assign label_5[150] = 10'b0000000001;
assign label_5[151] = 10'b0000000001;
assign label_5[152] = 10'b0000100000;
assign label_5[153] = 10'b0000000100;
assign label_5[154] = 10'b0000001000;
assign label_5[155] = 10'b0000001000;
assign label_5[156] = 10'b0000100000;
assign label_5[157] = 10'b0000001000;
assign label_5[158] = 10'b0000100000;
assign label_5[159] = 10'b0000000001;
assign label_5[160] = 10'b0000000001;
assign label_5[161] = 10'b0000000001;
assign label_5[162] = 10'b0000000100;
assign label_5[163] = 10'b0000010000;
assign label_5[164] = 10'b0000000001;
assign label_5[165] = 10'b0001000000;
assign label_5[166] = 10'b0000100000;
assign label_5[167] = 10'b0000000001;
assign label_5[168] = 10'b0000100000;
assign label_5[169] = 10'b0000000100;
assign label_5[170] = 10'b0000000001;
assign label_5[171] = 10'b0000000001;
assign label_5[172] = 10'b0000100000;
assign label_5[173] = 10'b0000000100;
assign label_5[174] = 10'b0000000001;
assign label_5[175] = 10'b0000001000;
assign label_5[176] = 10'b0000000001;
assign label_5[177] = 10'b0000000001;
assign label_5[178] = 10'b0001000000;
assign label_5[179] = 10'b0001000000;
assign label_5[180] = 10'b0000000001;
assign label_5[181] = 10'b0010000000;
assign label_5[182] = 10'b0000000001;
assign label_5[183] = 10'b0000000001;
assign label_5[184] = 10'b0000000001;
assign label_5[185] = 10'b0000000100;
assign label_5[186] = 10'b0000000001;
assign label_5[187] = 10'b0000000100;
assign label_5[188] = 10'b0000000001;
assign label_5[189] = 10'b0000000001;
assign label_5[190] = 10'b0000100000;
assign label_5[191] = 10'b0000000001;
assign label_5[192] = 10'b0000000100;
assign label_5[193] = 10'b0000000100;
assign label_5[194] = 10'b0010000000;
assign label_5[195] = 10'b0010000000;
assign label_5[196] = 10'b0000100000;
assign label_5[197] = 10'b0000000100;
assign label_5[198] = 10'b1000000000;
assign label_5[199] = 10'b0000000001;
assign label_5[200] = 10'b0000100000;
assign label_5[201] = 10'b0000000100;
assign label_5[202] = 10'b0000001000;
assign label_5[203] = 10'b0000100000;
assign label_5[204] = 10'b0000000100;
assign label_5[205] = 10'b0000000100;
assign label_5[206] = 10'b0000000100;
assign label_5[207] = 10'b0000000100;
assign label_5[208] = 10'b0000001000;
assign label_5[209] = 10'b0000100000;
assign label_5[210] = 10'b0000000001;
assign label_5[211] = 10'b0001000000;
assign label_5[212] = 10'b0001000000;
assign label_5[213] = 10'b0000000100;
assign label_5[214] = 10'b0000001000;
assign label_5[215] = 10'b0000000100;
assign label_5[216] = 10'b0000010000;
assign label_5[217] = 10'b0000010000;
assign label_5[218] = 10'b0000000001;
assign label_5[219] = 10'b0001000000;
assign label_5[220] = 10'b0000010000;
assign label_5[221] = 10'b0000000001;
assign label_5[222] = 10'b0000000001;
assign label_5[223] = 10'b0000000100;
assign label_5[224] = 10'b0000000100;
assign label_5[225] = 10'b0000000001;
assign label_5[226] = 10'b0000000100;
assign label_5[227] = 10'b0000010000;
assign label_5[228] = 10'b0000000001;
assign label_5[229] = 10'b0000000100;
assign label_5[230] = 10'b0000000001;
assign label_5[231] = 10'b0000000001;
assign label_5[232] = 10'b0000000100;
assign label_5[233] = 10'b0000000100;
assign label_5[234] = 10'b0000000001;
assign label_5[235] = 10'b0000000001;
assign label_5[236] = 10'b0000010000;
assign label_5[237] = 10'b0000010000;
assign label_5[238] = 10'b0000000001;
assign label_5[239] = 10'b0000000001;
assign label_5[240] = 10'b0001000000;
assign label_5[241] = 10'b0000000100;
assign label_5[242] = 10'b0000000001;
assign label_5[243] = 10'b0000000001;
assign label_5[244] = 10'b0000000001;
assign label_5[245] = 10'b0000000001;
assign label_5[246] = 10'b0000000100;
assign label_5[247] = 10'b0000000100;
assign label_5[248] = 10'b0000000001;
assign label_5[249] = 10'b0000000001;
assign label_5[250] = 10'b0000000100;
assign label_5[251] = 10'b0000001000;
assign label_5[252] = 10'b0000000100;
assign label_5[253] = 10'b0000000100;
assign label_5[254] = 10'b0000000100;
assign label_5[255] = 10'b0000000100;
assign label_5[256] = 10'b0000010000;
assign label_5[257] = 10'b0000010000;
assign label_5[258] = 10'b0000000100;
assign label_5[259] = 10'b0100000000;
assign label_5[260] = 10'b0000010000;
assign label_5[261] = 10'b1000000000;
assign label_5[262] = 10'b0000000100;
assign label_5[263] = 10'b0000010000;
assign label_5[264] = 10'b0000000100;
assign label_5[265] = 10'b0000000100;
assign label_5[266] = 10'b0001000000;
assign label_5[267] = 10'b0001000000;
assign label_5[268] = 10'b0000010000;
assign label_5[269] = 10'b0001000000;
assign label_5[270] = 10'b1000000000;
assign label_5[271] = 10'b0001000000;
assign label_5[272] = 10'b0000010000;
assign label_5[273] = 10'b0001000000;
assign label_5[274] = 10'b0000100000;
assign label_5[275] = 10'b1000000000;
assign label_5[276] = 10'b0001000000;
assign label_5[277] = 10'b0000100000;
assign label_5[278] = 10'b0001000000;
assign label_5[279] = 10'b0100000000;
assign label_5[280] = 10'b0000010000;
assign label_5[281] = 10'b0100000000;
assign label_5[282] = 10'b0000010000;
assign label_5[283] = 10'b0000010000;
assign label_5[284] = 10'b0100000000;
assign label_5[285] = 10'b0000010000;
assign label_5[286] = 10'b0000010000;
assign label_5[287] = 10'b0000000100;
assign label_5[288] = 10'b0001000000;
assign label_5[289] = 10'b0000010000;
assign label_5[290] = 10'b0001000000;
assign label_5[291] = 10'b0001000000;
assign label_5[292] = 10'b0001000000;
assign label_5[293] = 10'b0001000000;
assign label_5[294] = 10'b0000000010;
assign label_5[295] = 10'b0001000000;
assign label_5[296] = 10'b0001000000;
assign label_5[297] = 10'b0001000000;
assign label_5[298] = 10'b0001000000;
assign label_5[299] = 10'b0001000000;
assign label_5[300] = 10'b0000000100;
assign label_5[301] = 10'b0000000100;
assign label_5[302] = 10'b0000000100;
assign label_5[303] = 10'b0000000100;
assign label_5[304] = 10'b0000000100;
assign label_5[305] = 10'b0000000100;
assign label_5[306] = 10'b0000000100;
assign label_5[307] = 10'b0000000100;
assign label_5[308] = 10'b0000000100;
assign label_5[309] = 10'b0000000100;
assign label_5[310] = 10'b0000000100;
assign label_5[311] = 10'b0000000100;
assign label_5[312] = 10'b0000000100;
assign label_5[313] = 10'b0000000100;
assign label_5[314] = 10'b0000000100;
assign label_5[315] = 10'b0000000100;
assign label_5[316] = 10'b0000000100;
assign label_5[317] = 10'b0000000100;
assign label_5[318] = 10'b0000000100;
assign label_5[319] = 10'b0000000100;
assign label_5[320] = 10'b0001000000;
assign label_5[321] = 10'b0000100000;
assign label_5[322] = 10'b0001000000;
assign label_5[323] = 10'b0001000000;
assign label_5[324] = 10'b0001000000;
assign label_5[325] = 10'b0001000000;
assign label_5[326] = 10'b0001000000;
assign label_5[327] = 10'b0000100000;
assign label_5[328] = 10'b0000000100;
assign label_5[329] = 10'b0000000100;
assign label_5[330] = 10'b0000010000;
assign label_5[331] = 10'b0000010000;
assign label_5[332] = 10'b0001000000;
assign label_5[333] = 10'b0001000000;
assign label_5[334] = 10'b0001000000;
assign label_5[335] = 10'b0001000000;
assign label_5[336] = 10'b0000000100;
assign label_5[337] = 10'b0000000100;
assign label_5[338] = 10'b0000000100;
assign label_5[339] = 10'b0000000100;
assign label_5[340] = 10'b0001000000;
assign label_5[341] = 10'b0001000000;
assign label_5[342] = 10'b0000000100;
assign label_5[343] = 10'b0000000100;
assign label_5[344] = 10'b0001000000;
assign label_5[345] = 10'b0001000000;
assign label_5[346] = 10'b0000000100;
assign label_5[347] = 10'b0000000100;
assign label_5[348] = 10'b0000000001;
assign label_5[349] = 10'b0000000001;
assign label_5[350] = 10'b0001000000;
assign label_5[351] = 10'b0001000000;
assign label_5[352] = 10'b0000000100;
assign label_5[353] = 10'b0000000100;
assign label_5[354] = 10'b0000000100;
assign label_5[355] = 10'b0000000100;
assign label_5[356] = 10'b0000010000;
assign label_5[357] = 10'b0000010000;
assign label_5[358] = 10'b0000010000;
assign label_5[359] = 10'b0000010000;
assign label_5[360] = 10'b0000000100;
assign label_5[361] = 10'b0000000100;
assign label_5[362] = 10'b0000000100;
assign label_5[363] = 10'b0000000100;
assign label_5[364] = 10'b0000000100;
assign label_5[365] = 10'b0000000100;
assign label_5[366] = 10'b0000000100;
assign label_5[367] = 10'b0000000100;
assign label_5[368] = 10'b0001000000;
assign label_5[369] = 10'b0000010000;
assign label_5[370] = 10'b0001000000;
assign label_5[371] = 10'b0001000000;
assign label_5[372] = 10'b0000000100;
assign label_5[373] = 10'b0000000100;
assign label_5[374] = 10'b0000010000;
assign label_5[375] = 10'b0000010000;
assign label_5[376] = 10'b0000000100;
assign label_5[377] = 10'b0000000100;
assign label_5[378] = 10'b0000000100;
assign label_5[379] = 10'b0000000100;
assign label_5[380] = 10'b0001000000;
assign label_5[381] = 10'b0001000000;
assign label_5[382] = 10'b0000010000;
assign label_5[383] = 10'b0000000001;
assign label_5[384] = 10'b0010000000;
assign label_5[385] = 10'b0010000000;
assign label_5[386] = 10'b0000100000;
assign label_5[387] = 10'b0010000000;
assign label_5[388] = 10'b0000100000;
assign label_5[389] = 10'b0000000100;
assign label_5[390] = 10'b0001000000;
assign label_5[391] = 10'b0000000001;
assign label_5[392] = 10'b0000000100;
assign label_5[393] = 10'b0010000000;
assign label_5[394] = 10'b0000000010;
assign label_5[395] = 10'b0000000100;
assign label_5[396] = 10'b0000001000;
assign label_5[397] = 10'b0000000100;
assign label_5[398] = 10'b0000100000;
assign label_5[399] = 10'b0000000001;
assign label_5[400] = 10'b0010000000;
assign label_5[401] = 10'b1000000000;
assign label_5[402] = 10'b0010000000;
assign label_5[403] = 10'b1000000000;
assign label_5[404] = 10'b0001000000;
assign label_5[405] = 10'b0000000100;
assign label_5[406] = 10'b0000010000;
assign label_5[407] = 10'b1000000000;
assign label_5[408] = 10'b0000000100;
assign label_5[409] = 10'b0010000000;
assign label_5[410] = 10'b0100000000;
assign label_5[411] = 10'b0000100000;
assign label_5[412] = 10'b0000000001;
assign label_5[413] = 10'b1000000000;
assign label_5[414] = 10'b0001000000;
assign label_5[415] = 10'b0000000001;
assign label_5[416] = 10'b0000000100;
assign label_5[417] = 10'b0000000100;
assign label_5[418] = 10'b0010000000;
assign label_5[419] = 10'b0010000000;
assign label_5[420] = 10'b0000001000;
assign label_5[421] = 10'b1000000000;
assign label_5[422] = 10'b0000000100;
assign label_5[423] = 10'b0001000000;
assign label_5[424] = 10'b0000000001;
assign label_5[425] = 10'b0000000001;
assign label_5[426] = 10'b0000010000;
assign label_5[427] = 10'b0001000000;
assign label_5[428] = 10'b0000010000;
assign label_5[429] = 10'b1000000000;
assign label_5[430] = 10'b0000000100;
assign label_5[431] = 10'b0001000000;
assign label_5[432] = 10'b0010000000;
assign label_5[433] = 10'b1000000000;
assign label_5[434] = 10'b0100000000;
assign label_5[435] = 10'b0000000100;
assign label_5[436] = 10'b1000000000;
assign label_5[437] = 10'b0000000100;
assign label_5[438] = 10'b0000001000;
assign label_5[439] = 10'b0000010000;
assign label_5[440] = 10'b0000010000;
assign label_5[441] = 10'b1000000000;
assign label_5[442] = 10'b0010000000;
assign label_5[443] = 10'b1000000000;
assign label_5[444] = 10'b1000000000;
assign label_5[445] = 10'b1000000000;
assign label_5[446] = 10'b0000010000;
assign label_5[447] = 10'b1000000000;
assign label_5[448] = 10'b0000010000;
assign label_5[449] = 10'b0100000000;
assign label_5[450] = 10'b0000010000;
assign label_5[451] = 10'b0000010000;
assign label_5[452] = 10'b0000001000;
assign label_5[453] = 10'b0000100000;
assign label_5[454] = 10'b0100000000;
assign label_5[455] = 10'b0000010000;
assign label_5[456] = 10'b1000000000;
assign label_5[457] = 10'b0010000000;
assign label_5[458] = 10'b1000000000;
assign label_5[459] = 10'b1000000000;
assign label_5[460] = 10'b0000100000;
assign label_5[461] = 10'b0000001000;
assign label_5[462] = 10'b0000010000;
assign label_5[463] = 10'b1000000000;
assign label_5[464] = 10'b0000100000;
assign label_5[465] = 10'b0000010000;
assign label_5[466] = 10'b0000000100;
assign label_5[467] = 10'b0000001000;
assign label_5[468] = 10'b0000000100;
assign label_5[469] = 10'b0000000100;
assign label_5[470] = 10'b0000001000;
assign label_5[471] = 10'b0000100000;
assign label_5[472] = 10'b0000000001;
assign label_5[473] = 10'b0000000001;
assign label_5[474] = 10'b0000000100;
assign label_5[475] = 10'b0000000100;
assign label_5[476] = 10'b0000100000;
assign label_5[477] = 10'b0000001000;
assign label_5[478] = 10'b0100000000;
assign label_5[479] = 10'b0000000100;
assign label_5[480] = 10'b0000000100;
assign label_5[481] = 10'b0100000000;
assign label_5[482] = 10'b0000100000;
assign label_5[483] = 10'b0001000000;
assign label_5[484] = 10'b0000000100;
assign label_5[485] = 10'b0000001000;
assign label_5[486] = 10'b0000000100;
assign label_5[487] = 10'b0000000100;
assign label_5[488] = 10'b0000000100;
assign label_5[489] = 10'b0000100000;
assign label_5[490] = 10'b0100000000;
assign label_5[491] = 10'b0100000000;
assign label_5[492] = 10'b0000000100;
assign label_5[493] = 10'b0001000000;
assign label_5[494] = 10'b0000100000;
assign label_5[495] = 10'b0100000000;
assign label_5[496] = 10'b0000100000;
assign label_5[497] = 10'b0000000100;
assign label_5[498] = 10'b0100000000;
assign label_5[499] = 10'b0100000000;
assign label_5[500] = 10'b0000000100;
assign label_5[501] = 10'b0000010000;
assign label_5[502] = 10'b0000000100;
assign label_5[503] = 10'b0100000000;
assign label_5[504] = 10'b0000100000;
assign label_5[505] = 10'b0100000000;
assign label_5[506] = 10'b0000100000;
assign label_5[507] = 10'b0000000100;
assign label_5[508] = 10'b0000000001;
assign label_5[509] = 10'b0000000001;
assign label_5[510] = 10'b0000000100;
assign label_5[511] = 10'b0100000000;
assign label_5[512] = 10'b0000000010;
assign label_5[513] = 10'b0000001000;
assign label_5[514] = 10'b1000000000;
assign label_5[515] = 10'b0000001000;
assign label_5[516] = 10'b0000100000;
assign label_5[517] = 10'b0100000000;
assign label_5[518] = 10'b0000000100;
assign label_5[519] = 10'b0000001000;
assign label_5[520] = 10'b0000100000;
assign label_5[521] = 10'b0000001000;
assign label_5[522] = 10'b0000100000;
assign label_5[523] = 10'b1000000000;
assign label_5[524] = 10'b0000100000;
assign label_5[525] = 10'b0100000000;
assign label_5[526] = 10'b0100000000;
assign label_5[527] = 10'b0000000001;
assign label_5[528] = 10'b0000001000;
assign label_5[529] = 10'b0000000100;
assign label_5[530] = 10'b0000001000;
assign label_5[531] = 10'b0000001000;
assign label_5[532] = 10'b0000001000;
assign label_5[533] = 10'b1000000000;
assign label_5[534] = 10'b0000001000;
assign label_5[535] = 10'b0000001000;
assign label_5[536] = 10'b0000100000;
assign label_5[537] = 10'b0000100000;
assign label_5[538] = 10'b0000001000;
assign label_5[539] = 10'b0000100000;
assign label_5[540] = 10'b0000100000;
assign label_5[541] = 10'b0100000000;
assign label_5[542] = 10'b0000000001;
assign label_5[543] = 10'b0100000000;
assign label_5[544] = 10'b0000100000;
assign label_5[545] = 10'b0000001000;
assign label_5[546] = 10'b0000100000;
assign label_5[547] = 10'b0000100000;
assign label_5[548] = 10'b0000001000;
assign label_5[549] = 10'b1000000000;
assign label_5[550] = 10'b0000100000;
assign label_5[551] = 10'b0000000001;
assign label_5[552] = 10'b0000100000;
assign label_5[553] = 10'b1000000000;
assign label_5[554] = 10'b0000001000;
assign label_5[555] = 10'b0000100000;
assign label_5[556] = 10'b1000000000;
assign label_5[557] = 10'b1000000000;
assign label_5[558] = 10'b0000001000;
assign label_5[559] = 10'b0100000000;
assign label_5[560] = 10'b0000100000;
assign label_5[561] = 10'b0000100000;
assign label_5[562] = 10'b0000100000;
assign label_5[563] = 10'b1000000000;
assign label_5[564] = 10'b0000001000;
assign label_5[565] = 10'b0000100000;
assign label_5[566] = 10'b0000001000;
assign label_5[567] = 10'b0000001000;
assign label_5[568] = 10'b0000100000;
assign label_5[569] = 10'b0100000000;
assign label_5[570] = 10'b0000100000;
assign label_5[571] = 10'b0100000000;
assign label_5[572] = 10'b0100000000;
assign label_5[573] = 10'b0001000000;
assign label_5[574] = 10'b0000000001;
assign label_5[575] = 10'b0100000000;
assign label_5[576] = 10'b0000000010;
assign label_5[577] = 10'b0000100000;
assign label_5[578] = 10'b0000000100;
assign label_5[579] = 10'b0100000000;
assign label_5[580] = 10'b0000000100;
assign label_5[581] = 10'b0000010000;
assign label_5[582] = 10'b0100000000;
assign label_5[583] = 10'b0100000000;
assign label_5[584] = 10'b0001000000;
assign label_5[585] = 10'b0000100000;
assign label_5[586] = 10'b0000000100;
assign label_5[587] = 10'b0000001000;
assign label_5[588] = 10'b0000000100;
assign label_5[589] = 10'b0000001000;
assign label_5[590] = 10'b0100000000;
assign label_5[591] = 10'b0000000100;
assign label_5[592] = 10'b0000000010;
assign label_5[593] = 10'b0000001000;
assign label_5[594] = 10'b0000001000;
assign label_5[595] = 10'b0100000000;
assign label_5[596] = 10'b0000000100;
assign label_5[597] = 10'b0000001000;
assign label_5[598] = 10'b0000001000;
assign label_5[599] = 10'b0100000000;
assign label_5[600] = 10'b0100000000;
assign label_5[601] = 10'b0000100000;
assign label_5[602] = 10'b0100000000;
assign label_5[603] = 10'b0100000000;
assign label_5[604] = 10'b0001000000;
assign label_5[605] = 10'b0000100000;
assign label_5[606] = 10'b0000000100;
assign label_5[607] = 10'b0000001000;
assign label_5[608] = 10'b0000100000;
assign label_5[609] = 10'b0100000000;
assign label_5[610] = 10'b0001000000;
assign label_5[611] = 10'b0000100000;
assign label_5[612] = 10'b0000100000;
assign label_5[613] = 10'b0000100000;
assign label_5[614] = 10'b0001000000;
assign label_5[615] = 10'b0100000000;
assign label_5[616] = 10'b0001000000;
assign label_5[617] = 10'b0100000000;
assign label_5[618] = 10'b0000100000;
assign label_5[619] = 10'b0000000001;
assign label_5[620] = 10'b0100000000;
assign label_5[621] = 10'b0000000100;
assign label_5[622] = 10'b0100000000;
assign label_5[623] = 10'b0000001000;
assign label_5[624] = 10'b0000100000;
assign label_5[625] = 10'b0001000000;
assign label_5[626] = 10'b0001000000;
assign label_5[627] = 10'b0001000000;
assign label_5[628] = 10'b0100000000;
assign label_5[629] = 10'b0010000000;
assign label_5[630] = 10'b1000000000;
assign label_5[631] = 10'b0000000001;
assign label_5[632] = 10'b0000100000;
assign label_5[633] = 10'b0000000001;
assign label_5[634] = 10'b0001000000;
assign label_5[635] = 10'b0000000001;
assign label_5[636] = 10'b0000000001;
assign label_5[637] = 10'b0000001000;
assign label_5[638] = 10'b0000000001;
assign label_5[639] = 10'b0000000001;
assign label_5[640] = 10'b0000000010;
assign label_5[641] = 10'b0000000100;
assign label_5[642] = 10'b0000000010;
assign label_5[643] = 10'b0001000000;
assign label_5[644] = 10'b0000100000;
assign label_5[645] = 10'b0000000100;
assign label_5[646] = 10'b0000000100;
assign label_5[647] = 10'b0000000100;
assign label_5[648] = 10'b0100000000;
assign label_5[649] = 10'b1000000000;
assign label_5[650] = 10'b0100000000;
assign label_5[651] = 10'b0000001000;
assign label_5[652] = 10'b0000000010;
assign label_5[653] = 10'b0100000000;
assign label_5[654] = 10'b0000100000;
assign label_5[655] = 10'b0100000000;
assign label_5[656] = 10'b0010000000;
assign label_5[657] = 10'b0000000100;
assign label_5[658] = 10'b0010000000;
assign label_5[659] = 10'b0000001000;
assign label_5[660] = 10'b0010000000;
assign label_5[661] = 10'b0000000010;
assign label_5[662] = 10'b0100000000;
assign label_5[663] = 10'b0000001000;
assign label_5[664] = 10'b0000000100;
assign label_5[665] = 10'b1000000000;
assign label_5[666] = 10'b0000001000;
assign label_5[667] = 10'b0000000100;
assign label_5[668] = 10'b0001000000;
assign label_5[669] = 10'b0001000000;
assign label_5[670] = 10'b0001000000;
assign label_5[671] = 10'b0001000000;
assign label_5[672] = 10'b0000000010;
assign label_5[673] = 10'b0000000100;
assign label_5[674] = 10'b0100000000;
assign label_5[675] = 10'b0000000100;
assign label_5[676] = 10'b0000000100;
assign label_5[677] = 10'b0100000000;
assign label_5[678] = 10'b0000000100;
assign label_5[679] = 10'b0001000000;
assign label_5[680] = 10'b0000000100;
assign label_5[681] = 10'b0000000100;
assign label_5[682] = 10'b0000000100;
assign label_5[683] = 10'b0001000000;
assign label_5[684] = 10'b0100000000;
assign label_5[685] = 10'b0000001000;
assign label_5[686] = 10'b0000000100;
assign label_5[687] = 10'b0100000000;
assign label_5[688] = 10'b0000000100;
assign label_5[689] = 10'b0001000000;
assign label_5[690] = 10'b0001000000;
assign label_5[691] = 10'b0001000000;
assign label_5[692] = 10'b0001000000;
assign label_5[693] = 10'b0001000000;
assign label_5[694] = 10'b1000000000;
assign label_5[695] = 10'b1000000000;
assign label_5[696] = 10'b0001000000;
assign label_5[697] = 10'b0001000000;
assign label_5[698] = 10'b0001000000;
assign label_5[699] = 10'b0001000000;
assign label_5[700] = 10'b0000000001;
assign label_5[701] = 10'b0000000001;
assign label_5[702] = 10'b1000000000;
assign label_5[703] = 10'b1000000000;
assign label_5[704] = 10'b0000010000;
assign label_5[705] = 10'b0000100000;
assign label_5[706] = 10'b1000000000;
assign label_5[707] = 10'b0100000000;
assign label_5[708] = 10'b0000100000;
assign label_5[709] = 10'b0000100000;
assign label_5[710] = 10'b1000000000;
assign label_5[711] = 10'b0100000000;
assign label_5[712] = 10'b0000010000;
assign label_5[713] = 10'b0100000000;
assign label_5[714] = 10'b0001000000;
assign label_5[715] = 10'b0100000000;
assign label_5[716] = 10'b0100000000;
assign label_5[717] = 10'b0000000100;
assign label_5[718] = 10'b0100000000;
assign label_5[719] = 10'b0100000000;
assign label_5[720] = 10'b0000000010;
assign label_5[721] = 10'b0000010000;
assign label_5[722] = 10'b0000100000;
assign label_5[723] = 10'b0000100000;
assign label_5[724] = 10'b0100000000;
assign label_5[725] = 10'b0000100000;
assign label_5[726] = 10'b0100000000;
assign label_5[727] = 10'b0001000000;
assign label_5[728] = 10'b0100000000;
assign label_5[729] = 10'b0100000000;
assign label_5[730] = 10'b0000000100;
assign label_5[731] = 10'b0000100000;
assign label_5[732] = 10'b0000000001;
assign label_5[733] = 10'b0000000100;
assign label_5[734] = 10'b0000000010;
assign label_5[735] = 10'b0100000000;
assign label_5[736] = 10'b0000010000;
assign label_5[737] = 10'b0001000000;
assign label_5[738] = 10'b0001000000;
assign label_5[739] = 10'b0001000000;
assign label_5[740] = 10'b0000000100;
assign label_5[741] = 10'b0000000100;
assign label_5[742] = 10'b0000000001;
assign label_5[743] = 10'b0001000000;
assign label_5[744] = 10'b1000000000;
assign label_5[745] = 10'b0000010000;
assign label_5[746] = 10'b0000000100;
assign label_5[747] = 10'b0010000000;
assign label_5[748] = 10'b0000010000;
assign label_5[749] = 10'b0000000100;
assign label_5[750] = 10'b0000010000;
assign label_5[751] = 10'b0001000000;
assign label_5[752] = 10'b0001000000;
assign label_5[753] = 10'b1000000000;
assign label_5[754] = 10'b0000100000;
assign label_5[755] = 10'b0001000000;
assign label_5[756] = 10'b0001000000;
assign label_5[757] = 10'b0000010000;
assign label_5[758] = 10'b0001000000;
assign label_5[759] = 10'b0000000001;
assign label_5[760] = 10'b0000100000;
assign label_5[761] = 10'b0000100000;
assign label_5[762] = 10'b0000010000;
assign label_5[763] = 10'b0000000100;
assign label_5[764] = 10'b0000000001;
assign label_5[765] = 10'b0000000100;
assign label_5[766] = 10'b0000000001;
assign label_5[767] = 10'b0000000001;
assign label_5[768] = 10'b0010000000;
assign label_5[769] = 10'b0000010000;
assign label_5[770] = 10'b0000010000;
assign label_5[771] = 10'b0010000000;
assign label_5[772] = 10'b0000010000;
assign label_5[773] = 10'b0000100000;
assign label_5[774] = 10'b0010000000;
assign label_5[775] = 10'b0000010000;
assign label_5[776] = 10'b0000100000;
assign label_5[777] = 10'b0100000000;
assign label_5[778] = 10'b0000010000;
assign label_5[779] = 10'b1000000000;
assign label_5[780] = 10'b0000001000;
assign label_5[781] = 10'b0000100000;
assign label_5[782] = 10'b1000000000;
assign label_5[783] = 10'b0010000000;
assign label_5[784] = 10'b1000000000;
assign label_5[785] = 10'b0000100000;
assign label_5[786] = 10'b1000000000;
assign label_5[787] = 10'b0010000000;
assign label_5[788] = 10'b1000000000;
assign label_5[789] = 10'b0000010000;
assign label_5[790] = 10'b0000100000;
assign label_5[791] = 10'b0000001000;
assign label_5[792] = 10'b0000100000;
assign label_5[793] = 10'b0000001000;
assign label_5[794] = 10'b0001000000;
assign label_5[795] = 10'b0001000000;
assign label_5[796] = 10'b0000001000;
assign label_5[797] = 10'b0000001000;
assign label_5[798] = 10'b0000000100;
assign label_5[799] = 10'b0000001000;
assign label_5[800] = 10'b0000100000;
assign label_5[801] = 10'b0000100000;
assign label_5[802] = 10'b0000001000;
assign label_5[803] = 10'b0000100000;
assign label_5[804] = 10'b0000001000;
assign label_5[805] = 10'b0000100000;
assign label_5[806] = 10'b0001000000;
assign label_5[807] = 10'b0000001000;
assign label_5[808] = 10'b0000001000;
assign label_5[809] = 10'b0000000100;
assign label_5[810] = 10'b0000001000;
assign label_5[811] = 10'b0000001000;
assign label_5[812] = 10'b0000000100;
assign label_5[813] = 10'b0000000100;
assign label_5[814] = 10'b0000000100;
assign label_5[815] = 10'b0000000100;
assign label_5[816] = 10'b0000001000;
assign label_5[817] = 10'b0000100000;
assign label_5[818] = 10'b0000000001;
assign label_5[819] = 10'b0000000001;
assign label_5[820] = 10'b0000000001;
assign label_5[821] = 10'b0000001000;
assign label_5[822] = 10'b0000001000;
assign label_5[823] = 10'b0000000100;
assign label_5[824] = 10'b0000100000;
assign label_5[825] = 10'b0000100000;
assign label_5[826] = 10'b0000100000;
assign label_5[827] = 10'b0000000001;
assign label_5[828] = 10'b0000001000;
assign label_5[829] = 10'b0000001000;
assign label_5[830] = 10'b0000000100;
assign label_5[831] = 10'b0000000100;
assign label_5[832] = 10'b0000100000;
assign label_5[833] = 10'b0000001000;
assign label_5[834] = 10'b0000000100;
assign label_5[835] = 10'b0001000000;
assign label_5[836] = 10'b0000100000;
assign label_5[837] = 10'b0000001000;
assign label_5[838] = 10'b1000000000;
assign label_5[839] = 10'b0001000000;
assign label_5[840] = 10'b0000100000;
assign label_5[841] = 10'b0000000100;
assign label_5[842] = 10'b0000100000;
assign label_5[843] = 10'b0000100000;
assign label_5[844] = 10'b0000100000;
assign label_5[845] = 10'b0000001000;
assign label_5[846] = 10'b0000100000;
assign label_5[847] = 10'b0000100000;
assign label_5[848] = 10'b0000001000;
assign label_5[849] = 10'b0000001000;
assign label_5[850] = 10'b0100000000;
assign label_5[851] = 10'b0000001000;
assign label_5[852] = 10'b0000000100;
assign label_5[853] = 10'b0000000100;
assign label_5[854] = 10'b0000000100;
assign label_5[855] = 10'b0000000100;
assign label_5[856] = 10'b0000001000;
assign label_5[857] = 10'b0000000100;
assign label_5[858] = 10'b0000010000;
assign label_5[859] = 10'b0000000100;
assign label_5[860] = 10'b0000010000;
assign label_5[861] = 10'b0100000000;
assign label_5[862] = 10'b0000001000;
assign label_5[863] = 10'b0100000000;
assign label_5[864] = 10'b0000001000;
assign label_5[865] = 10'b0000010000;
assign label_5[866] = 10'b1000000000;
assign label_5[867] = 10'b0000000100;
assign label_5[868] = 10'b1000000000;
assign label_5[869] = 10'b0000100000;
assign label_5[870] = 10'b0000000100;
assign label_5[871] = 10'b0000001000;
assign label_5[872] = 10'b0000000100;
assign label_5[873] = 10'b0000000100;
assign label_5[874] = 10'b0000000100;
assign label_5[875] = 10'b0000000100;
assign label_5[876] = 10'b0000000100;
assign label_5[877] = 10'b0000000100;
assign label_5[878] = 10'b0000000100;
assign label_5[879] = 10'b0000000100;
assign label_5[880] = 10'b0000100000;
assign label_5[881] = 10'b0000001000;
assign label_5[882] = 10'b0100000000;
assign label_5[883] = 10'b0000001000;
assign label_5[884] = 10'b0000001000;
assign label_5[885] = 10'b0100000000;
assign label_5[886] = 10'b0000100000;
assign label_5[887] = 10'b0000100000;
assign label_5[888] = 10'b0000001000;
assign label_5[889] = 10'b0000001000;
assign label_5[890] = 10'b0000000100;
assign label_5[891] = 10'b0000001000;
assign label_5[892] = 10'b0000100000;
assign label_5[893] = 10'b0000100000;
assign label_5[894] = 10'b0000001000;
assign label_5[895] = 10'b0000100000;
assign label_5[896] = 10'b0000010000;
assign label_5[897] = 10'b1000000000;
assign label_5[898] = 10'b0001000000;
assign label_5[899] = 10'b0000010000;
assign label_5[900] = 10'b0001000000;
assign label_5[901] = 10'b0001000000;
assign label_5[902] = 10'b0001000000;
assign label_5[903] = 10'b0000000100;
assign label_5[904] = 10'b0001000000;
assign label_5[905] = 10'b0000010000;
assign label_5[906] = 10'b0001000000;
assign label_5[907] = 10'b0100000000;
assign label_5[908] = 10'b0001000000;
assign label_5[909] = 10'b0001000000;
assign label_5[910] = 10'b0001000000;
assign label_5[911] = 10'b0000000100;
assign label_5[912] = 10'b0000010000;
assign label_5[913] = 10'b0000010000;
assign label_5[914] = 10'b0000010000;
assign label_5[915] = 10'b0010000000;
assign label_5[916] = 10'b0010000000;
assign label_5[917] = 10'b0000010000;
assign label_5[918] = 10'b1000000000;
assign label_5[919] = 10'b0001000000;
assign label_5[920] = 10'b0000100000;
assign label_5[921] = 10'b0100000000;
assign label_5[922] = 10'b0000001000;
assign label_5[923] = 10'b0000100000;
assign label_5[924] = 10'b0100000000;
assign label_5[925] = 10'b0000100000;
assign label_5[926] = 10'b0100000000;
assign label_5[927] = 10'b0000001000;
assign label_5[928] = 10'b0000010000;
assign label_5[929] = 10'b0001000000;
assign label_5[930] = 10'b0000010000;
assign label_5[931] = 10'b1000000000;
assign label_5[932] = 10'b0000000100;
assign label_5[933] = 10'b0000000100;
assign label_5[934] = 10'b0000010000;
assign label_5[935] = 10'b0000000001;
assign label_5[936] = 10'b1000000000;
assign label_5[937] = 10'b1000000000;
assign label_5[938] = 10'b0000010000;
assign label_5[939] = 10'b1000000000;
assign label_5[940] = 10'b0000000100;
assign label_5[941] = 10'b1000000000;
assign label_5[942] = 10'b1000000000;
assign label_5[943] = 10'b0000010000;
assign label_5[944] = 10'b0100000000;
assign label_5[945] = 10'b0100000000;
assign label_5[946] = 10'b0000000100;
assign label_5[947] = 10'b0000000100;
assign label_5[948] = 10'b0001000000;
assign label_5[949] = 10'b0100000000;
assign label_5[950] = 10'b0100000000;
assign label_5[951] = 10'b0100000000;
assign label_5[952] = 10'b0000000100;
assign label_5[953] = 10'b0000000100;
assign label_5[954] = 10'b0000001000;
assign label_5[955] = 10'b0000000100;
assign label_5[956] = 10'b0000000100;
assign label_5[957] = 10'b0000010000;
assign label_5[958] = 10'b0100000000;
assign label_5[959] = 10'b0001000000;
assign label_5[960] = 10'b0100000000;
assign label_5[961] = 10'b0000000010;
assign label_5[962] = 10'b0100000000;
assign label_5[963] = 10'b0100000000;
assign label_5[964] = 10'b0000001000;
assign label_5[965] = 10'b0000100000;
assign label_5[966] = 10'b0000001000;
assign label_5[967] = 10'b0100000000;
assign label_5[968] = 10'b0010000000;
assign label_5[969] = 10'b0000001000;
assign label_5[970] = 10'b0100000000;
assign label_5[971] = 10'b0000001000;
assign label_5[972] = 10'b0000001000;
assign label_5[973] = 10'b0000000100;
assign label_5[974] = 10'b0000000100;
assign label_5[975] = 10'b0000001000;
assign label_5[976] = 10'b1000000000;
assign label_5[977] = 10'b0100000000;
assign label_5[978] = 10'b0100000000;
assign label_5[979] = 10'b0100000000;
assign label_5[980] = 10'b0100000000;
assign label_5[981] = 10'b0100000000;
assign label_5[982] = 10'b0100000000;
assign label_5[983] = 10'b0000001000;
assign label_5[984] = 10'b0100000000;
assign label_5[985] = 10'b0000100000;
assign label_5[986] = 10'b0100000000;
assign label_5[987] = 10'b0100000000;
assign label_5[988] = 10'b0100000000;
assign label_5[989] = 10'b0100000000;
assign label_5[990] = 10'b0001000000;
assign label_5[991] = 10'b0001000000;
assign label_5[992] = 10'b1000000000;
assign label_5[993] = 10'b0000010000;
assign label_5[994] = 10'b0100000000;
assign label_5[995] = 10'b1000000000;
assign label_5[996] = 10'b0000001000;
assign label_5[997] = 10'b1000000000;
assign label_5[998] = 10'b0000100000;
assign label_5[999] = 10'b0100000000;
assign label_5[1000] = 10'b0000000001;
assign label_5[1001] = 10'b0000000001;
assign label_5[1002] = 10'b0000000001;
assign label_5[1003] = 10'b0000000001;
assign label_5[1004] = 10'b0000000100;
assign label_5[1005] = 10'b0000000100;
assign label_5[1006] = 10'b0100000000;
assign label_5[1007] = 10'b0000000100;
assign label_5[1008] = 10'b0000010000;
assign label_5[1009] = 10'b0000001000;
assign label_5[1010] = 10'b0000000001;
assign label_5[1011] = 10'b0000000001;
assign label_5[1012] = 10'b0100000000;
assign label_5[1013] = 10'b0100000000;
assign label_5[1014] = 10'b0000001000;
assign label_5[1015] = 10'b0000001000;
assign label_5[1016] = 10'b0000010000;
assign label_5[1017] = 10'b0100000000;
assign label_5[1018] = 10'b0000001000;
assign label_5[1019] = 10'b0000000001;
assign label_5[1020] = 10'b0000010000;
assign label_5[1021] = 10'b0000001000;
assign label_5[1022] = 10'b0100000000;
assign label_5[1023] = 10'b0000000001;
assign label_6[0] = 10'b0000100000;
assign label_6[1] = 10'b0000000100;
assign label_6[2] = 10'b0001000000;
assign label_6[3] = 10'b0000000100;
assign label_6[4] = 10'b0000000010;
assign label_6[5] = 10'b0000000100;
assign label_6[6] = 10'b0000000010;
assign label_6[7] = 10'b0000000100;
assign label_6[8] = 10'b0010000000;
assign label_6[9] = 10'b0000000100;
assign label_6[10] = 10'b0000000100;
assign label_6[11] = 10'b0000001000;
assign label_6[12] = 10'b1000000000;
assign label_6[13] = 10'b0000000001;
assign label_6[14] = 10'b0000010000;
assign label_6[15] = 10'b0000010000;
assign label_6[16] = 10'b0000000010;
assign label_6[17] = 10'b0001000000;
assign label_6[18] = 10'b0000000010;
assign label_6[19] = 10'b0100000000;
assign label_6[20] = 10'b0000000100;
assign label_6[21] = 10'b1000000000;
assign label_6[22] = 10'b0000001000;
assign label_6[23] = 10'b0000001000;
assign label_6[24] = 10'b0010000000;
assign label_6[25] = 10'b0100000000;
assign label_6[26] = 10'b0000001000;
assign label_6[27] = 10'b0000000100;
assign label_6[28] = 10'b0000000100;
assign label_6[29] = 10'b0010000000;
assign label_6[30] = 10'b0010000000;
assign label_6[31] = 10'b0100000000;
assign label_6[32] = 10'b0000000010;
assign label_6[33] = 10'b0000001000;
assign label_6[34] = 10'b0000001000;
assign label_6[35] = 10'b0000001000;
assign label_6[36] = 10'b0000001000;
assign label_6[37] = 10'b0000001000;
assign label_6[38] = 10'b0001000000;
assign label_6[39] = 10'b0000000001;
assign label_6[40] = 10'b0000100000;
assign label_6[41] = 10'b1000000000;
assign label_6[42] = 10'b0000000001;
assign label_6[43] = 10'b0100000000;
assign label_6[44] = 10'b0010000000;
assign label_6[45] = 10'b0000100000;
assign label_6[46] = 10'b0000000001;
assign label_6[47] = 10'b0000100000;
assign label_6[48] = 10'b0000000100;
assign label_6[49] = 10'b0000100000;
assign label_6[50] = 10'b0000001000;
assign label_6[51] = 10'b0100000000;
assign label_6[52] = 10'b0000000100;
assign label_6[53] = 10'b0001000000;
assign label_6[54] = 10'b0001000000;
assign label_6[55] = 10'b0000000100;
assign label_6[56] = 10'b0000000010;
assign label_6[57] = 10'b0100000000;
assign label_6[58] = 10'b0000000100;
assign label_6[59] = 10'b0000000100;
assign label_6[60] = 10'b0000000100;
assign label_6[61] = 10'b0000000100;
assign label_6[62] = 10'b0000000100;
assign label_6[63] = 10'b0000000100;
assign label_6[64] = 10'b0000010000;
assign label_6[65] = 10'b0000000100;
assign label_6[66] = 10'b0001000000;
assign label_6[67] = 10'b0000000010;
assign label_6[68] = 10'b0000010000;
assign label_6[69] = 10'b0000001000;
assign label_6[70] = 10'b0000000100;
assign label_6[71] = 10'b0001000000;
assign label_6[72] = 10'b0000000100;
assign label_6[73] = 10'b0000000100;
assign label_6[74] = 10'b0000010000;
assign label_6[75] = 10'b0000000010;
assign label_6[76] = 10'b0000001000;
assign label_6[77] = 10'b0001000000;
assign label_6[78] = 10'b0001000000;
assign label_6[79] = 10'b0000000010;
assign label_6[80] = 10'b0000000010;
assign label_6[81] = 10'b1000000000;
assign label_6[82] = 10'b0001000000;
assign label_6[83] = 10'b0100000000;
assign label_6[84] = 10'b0000010000;
assign label_6[85] = 10'b0100000000;
assign label_6[86] = 10'b0000001000;
assign label_6[87] = 10'b0000000100;
assign label_6[88] = 10'b0010000000;
assign label_6[89] = 10'b0000001000;
assign label_6[90] = 10'b0000000100;
assign label_6[91] = 10'b0000000100;
assign label_6[92] = 10'b0100000000;
assign label_6[93] = 10'b0000100000;
assign label_6[94] = 10'b0000001000;
assign label_6[95] = 10'b0000001000;
assign label_6[96] = 10'b0010000000;
assign label_6[97] = 10'b0010000000;
assign label_6[98] = 10'b0000001000;
assign label_6[99] = 10'b0000000100;
assign label_6[100] = 10'b0000010000;
assign label_6[101] = 10'b0000010000;
assign label_6[102] = 10'b0000000100;
assign label_6[103] = 10'b1000000000;
assign label_6[104] = 10'b0010000000;
assign label_6[105] = 10'b0000000100;
assign label_6[106] = 10'b0000001000;
assign label_6[107] = 10'b0000001000;
assign label_6[108] = 10'b1000000000;
assign label_6[109] = 10'b0000010000;
assign label_6[110] = 10'b0000001000;
assign label_6[111] = 10'b0100000000;
assign label_6[112] = 10'b0000001000;
assign label_6[113] = 10'b0000100000;
assign label_6[114] = 10'b0000010000;
assign label_6[115] = 10'b0000000001;
assign label_6[116] = 10'b0000000100;
assign label_6[117] = 10'b0000000100;
assign label_6[118] = 10'b0000000010;
assign label_6[119] = 10'b0000001000;
assign label_6[120] = 10'b0000000100;
assign label_6[121] = 10'b0000000100;
assign label_6[122] = 10'b0000001000;
assign label_6[123] = 10'b0100000000;
assign label_6[124] = 10'b0000001000;
assign label_6[125] = 10'b0100000000;
assign label_6[126] = 10'b0100000000;
assign label_6[127] = 10'b0000001000;
assign label_6[128] = 10'b0000100000;
assign label_6[129] = 10'b0000010000;
assign label_6[130] = 10'b0000010000;
assign label_6[131] = 10'b0001000000;
assign label_6[132] = 10'b0000010000;
assign label_6[133] = 10'b1000000000;
assign label_6[134] = 10'b0000010000;
assign label_6[135] = 10'b0000010000;
assign label_6[136] = 10'b0000100000;
assign label_6[137] = 10'b0000001000;
assign label_6[138] = 10'b0000100000;
assign label_6[139] = 10'b0000001000;
assign label_6[140] = 10'b0000001000;
assign label_6[141] = 10'b0000100000;
assign label_6[142] = 10'b0000010000;
assign label_6[143] = 10'b0100000000;
assign label_6[144] = 10'b0000010000;
assign label_6[145] = 10'b0001000000;
assign label_6[146] = 10'b0001000000;
assign label_6[147] = 10'b0001000000;
assign label_6[148] = 10'b0000000001;
assign label_6[149] = 10'b0000001000;
assign label_6[150] = 10'b0001000000;
assign label_6[151] = 10'b0100000000;
assign label_6[152] = 10'b0000001000;
assign label_6[153] = 10'b0001000000;
assign label_6[154] = 10'b0000100000;
assign label_6[155] = 10'b0000000100;
assign label_6[156] = 10'b0000000100;
assign label_6[157] = 10'b0000000001;
assign label_6[158] = 10'b0000100000;
assign label_6[159] = 10'b0000000100;
assign label_6[160] = 10'b0000001000;
assign label_6[161] = 10'b0000000100;
assign label_6[162] = 10'b0100000000;
assign label_6[163] = 10'b0000100000;
assign label_6[164] = 10'b0000001000;
assign label_6[165] = 10'b0000100000;
assign label_6[166] = 10'b0000001000;
assign label_6[167] = 10'b0100000000;
assign label_6[168] = 10'b0000010000;
assign label_6[169] = 10'b0100000000;
assign label_6[170] = 10'b0000001000;
assign label_6[171] = 10'b0100000000;
assign label_6[172] = 10'b0001000000;
assign label_6[173] = 10'b0001000000;
assign label_6[174] = 10'b0001000000;
assign label_6[175] = 10'b0001000000;
assign label_6[176] = 10'b0000001000;
assign label_6[177] = 10'b0000100000;
assign label_6[178] = 10'b0000001000;
assign label_6[179] = 10'b0000001000;
assign label_6[180] = 10'b0000001000;
assign label_6[181] = 10'b0000001000;
assign label_6[182] = 10'b0000001000;
assign label_6[183] = 10'b0100000000;
assign label_6[184] = 10'b0000001000;
assign label_6[185] = 10'b0000100000;
assign label_6[186] = 10'b0000100000;
assign label_6[187] = 10'b0100000000;
assign label_6[188] = 10'b0000001000;
assign label_6[189] = 10'b0000000100;
assign label_6[190] = 10'b0100000000;
assign label_6[191] = 10'b0000001000;
assign label_6[192] = 10'b1000000000;
assign label_6[193] = 10'b0000010000;
assign label_6[194] = 10'b0010000000;
assign label_6[195] = 10'b0000001000;
assign label_6[196] = 10'b1000000000;
assign label_6[197] = 10'b0000010000;
assign label_6[198] = 10'b0000001000;
assign label_6[199] = 10'b0000001000;
assign label_6[200] = 10'b0010000000;
assign label_6[201] = 10'b0000100000;
assign label_6[202] = 10'b0000010000;
assign label_6[203] = 10'b0000010000;
assign label_6[204] = 10'b0000010000;
assign label_6[205] = 10'b0000010000;
assign label_6[206] = 10'b0000010000;
assign label_6[207] = 10'b0000010000;
assign label_6[208] = 10'b0010000000;
assign label_6[209] = 10'b0010000000;
assign label_6[210] = 10'b0000100000;
assign label_6[211] = 10'b0000100000;
assign label_6[212] = 10'b0000010000;
assign label_6[213] = 10'b0000010000;
assign label_6[214] = 10'b0010000000;
assign label_6[215] = 10'b0010000000;
assign label_6[216] = 10'b0000010000;
assign label_6[217] = 10'b0000010000;
assign label_6[218] = 10'b0000010000;
assign label_6[219] = 10'b0000010000;
assign label_6[220] = 10'b0000100000;
assign label_6[221] = 10'b0000100000;
assign label_6[222] = 10'b0000100000;
assign label_6[223] = 10'b0000100000;
assign label_6[224] = 10'b0000100000;
assign label_6[225] = 10'b0000001000;
assign label_6[226] = 10'b0000100000;
assign label_6[227] = 10'b0010000000;
assign label_6[228] = 10'b0010000000;
assign label_6[229] = 10'b0000100000;
assign label_6[230] = 10'b0010000000;
assign label_6[231] = 10'b0100000000;
assign label_6[232] = 10'b0000001000;
assign label_6[233] = 10'b0000001000;
assign label_6[234] = 10'b0000001000;
assign label_6[235] = 10'b0000001000;
assign label_6[236] = 10'b0000001000;
assign label_6[237] = 10'b0000001000;
assign label_6[238] = 10'b0000001000;
assign label_6[239] = 10'b0000001000;
assign label_6[240] = 10'b0000001000;
assign label_6[241] = 10'b0000001000;
assign label_6[242] = 10'b0010000000;
assign label_6[243] = 10'b0100000000;
assign label_6[244] = 10'b0100000000;
assign label_6[245] = 10'b1000000000;
assign label_6[246] = 10'b0000100000;
assign label_6[247] = 10'b0100000000;
assign label_6[248] = 10'b0010000000;
assign label_6[249] = 10'b1000000000;
assign label_6[250] = 10'b0010000000;
assign label_6[251] = 10'b1000000000;
assign label_6[252] = 10'b1000000000;
assign label_6[253] = 10'b0100000000;
assign label_6[254] = 10'b1000000000;
assign label_6[255] = 10'b0000100000;
assign label_6[256] = 10'b0010000000;
assign label_6[257] = 10'b0000000100;
assign label_6[258] = 10'b0010000000;
assign label_6[259] = 10'b0000000001;
assign label_6[260] = 10'b1000000000;
assign label_6[261] = 10'b0001000000;
assign label_6[262] = 10'b1000000000;
assign label_6[263] = 10'b0000000001;
assign label_6[264] = 10'b0010000000;
assign label_6[265] = 10'b0000001000;
assign label_6[266] = 10'b0000100000;
assign label_6[267] = 10'b0000001000;
assign label_6[268] = 10'b0000100000;
assign label_6[269] = 10'b0100000000;
assign label_6[270] = 10'b1000000000;
assign label_6[271] = 10'b0010000000;
assign label_6[272] = 10'b0000001000;
assign label_6[273] = 10'b0000000001;
assign label_6[274] = 10'b0000000100;
assign label_6[275] = 10'b0001000000;
assign label_6[276] = 10'b0000000001;
assign label_6[277] = 10'b0000000001;
assign label_6[278] = 10'b0000000001;
assign label_6[279] = 10'b0000000100;
assign label_6[280] = 10'b0000100000;
assign label_6[281] = 10'b0100000000;
assign label_6[282] = 10'b0000000001;
assign label_6[283] = 10'b0000000001;
assign label_6[284] = 10'b0100000000;
assign label_6[285] = 10'b0100000000;
assign label_6[286] = 10'b0100000000;
assign label_6[287] = 10'b0100000000;
assign label_6[288] = 10'b0000000001;
assign label_6[289] = 10'b0000100000;
assign label_6[290] = 10'b0000000100;
assign label_6[291] = 10'b0001000000;
assign label_6[292] = 10'b0001000000;
assign label_6[293] = 10'b0000000100;
assign label_6[294] = 10'b0000000100;
assign label_6[295] = 10'b0100000000;
assign label_6[296] = 10'b0000100000;
assign label_6[297] = 10'b0000001000;
assign label_6[298] = 10'b0100000000;
assign label_6[299] = 10'b0000010000;
assign label_6[300] = 10'b0000001000;
assign label_6[301] = 10'b0000100000;
assign label_6[302] = 10'b0100000000;
assign label_6[303] = 10'b0000000001;
assign label_6[304] = 10'b0000100000;
assign label_6[305] = 10'b0000001000;
assign label_6[306] = 10'b0000100000;
assign label_6[307] = 10'b0000001000;
assign label_6[308] = 10'b0000100000;
assign label_6[309] = 10'b0000001000;
assign label_6[310] = 10'b0000001000;
assign label_6[311] = 10'b0000001000;
assign label_6[312] = 10'b0000000100;
assign label_6[313] = 10'b0001000000;
assign label_6[314] = 10'b0001000000;
assign label_6[315] = 10'b0000010000;
assign label_6[316] = 10'b0100000000;
assign label_6[317] = 10'b0000001000;
assign label_6[318] = 10'b0100000000;
assign label_6[319] = 10'b0000100000;
assign label_6[320] = 10'b0000010000;
assign label_6[321] = 10'b0000010000;
assign label_6[322] = 10'b0001000000;
assign label_6[323] = 10'b0000100000;
assign label_6[324] = 10'b0000010000;
assign label_6[325] = 10'b1000000000;
assign label_6[326] = 10'b1000000000;
assign label_6[327] = 10'b0100000000;
assign label_6[328] = 10'b0000010000;
assign label_6[329] = 10'b0000000001;
assign label_6[330] = 10'b0000001000;
assign label_6[331] = 10'b0000100000;
assign label_6[332] = 10'b0000010000;
assign label_6[333] = 10'b0100000000;
assign label_6[334] = 10'b0100000000;
assign label_6[335] = 10'b0000010000;
assign label_6[336] = 10'b0000010000;
assign label_6[337] = 10'b0000100000;
assign label_6[338] = 10'b0001000000;
assign label_6[339] = 10'b0001000000;
assign label_6[340] = 10'b0000000001;
assign label_6[341] = 10'b0000100000;
assign label_6[342] = 10'b0100000000;
assign label_6[343] = 10'b0100000000;
assign label_6[344] = 10'b0000100000;
assign label_6[345] = 10'b0000100000;
assign label_6[346] = 10'b0000100000;
assign label_6[347] = 10'b0100000000;
assign label_6[348] = 10'b0010000000;
assign label_6[349] = 10'b0010000000;
assign label_6[350] = 10'b0000010000;
assign label_6[351] = 10'b0000100000;
assign label_6[352] = 10'b0000010000;
assign label_6[353] = 10'b0100000000;
assign label_6[354] = 10'b0000001000;
assign label_6[355] = 10'b0000100000;
assign label_6[356] = 10'b1000000000;
assign label_6[357] = 10'b0010000000;
assign label_6[358] = 10'b0000100000;
assign label_6[359] = 10'b1000000000;
assign label_6[360] = 10'b0000001000;
assign label_6[361] = 10'b0000100000;
assign label_6[362] = 10'b0100000000;
assign label_6[363] = 10'b0100000000;
assign label_6[364] = 10'b0000100000;
assign label_6[365] = 10'b0000001000;
assign label_6[366] = 10'b0000000100;
assign label_6[367] = 10'b0000000001;
assign label_6[368] = 10'b1000000000;
assign label_6[369] = 10'b0000001000;
assign label_6[370] = 10'b0000000001;
assign label_6[371] = 10'b1000000000;
assign label_6[372] = 10'b0100000000;
assign label_6[373] = 10'b0000010000;
assign label_6[374] = 10'b0100000000;
assign label_6[375] = 10'b0000001000;
assign label_6[376] = 10'b0000100000;
assign label_6[377] = 10'b0000001000;
assign label_6[378] = 10'b0100000000;
assign label_6[379] = 10'b0000100000;
assign label_6[380] = 10'b0010000000;
assign label_6[381] = 10'b0000000001;
assign label_6[382] = 10'b0100000000;
assign label_6[383] = 10'b0000001000;
assign label_6[384] = 10'b0000010000;
assign label_6[385] = 10'b0000010000;
assign label_6[386] = 10'b0001000000;
assign label_6[387] = 10'b0000010000;
assign label_6[388] = 10'b0000100000;
assign label_6[389] = 10'b0100000000;
assign label_6[390] = 10'b0100000000;
assign label_6[391] = 10'b0000001000;
assign label_6[392] = 10'b0000010000;
assign label_6[393] = 10'b0000100000;
assign label_6[394] = 10'b0001000000;
assign label_6[395] = 10'b0000010000;
assign label_6[396] = 10'b1000000000;
assign label_6[397] = 10'b0000010000;
assign label_6[398] = 10'b0001000000;
assign label_6[399] = 10'b0001000000;
assign label_6[400] = 10'b0100000000;
assign label_6[401] = 10'b0000100000;
assign label_6[402] = 10'b0000000100;
assign label_6[403] = 10'b0100000000;
assign label_6[404] = 10'b0100000000;
assign label_6[405] = 10'b0100000000;
assign label_6[406] = 10'b0010000000;
assign label_6[407] = 10'b0010000000;
assign label_6[408] = 10'b0000010000;
assign label_6[409] = 10'b0000001000;
assign label_6[410] = 10'b0100000000;
assign label_6[411] = 10'b0100000000;
assign label_6[412] = 10'b0001000000;
assign label_6[413] = 10'b0000010000;
assign label_6[414] = 10'b0100000000;
assign label_6[415] = 10'b0000010000;
assign label_6[416] = 10'b0001000000;
assign label_6[417] = 10'b0000100000;
assign label_6[418] = 10'b0000000001;
assign label_6[419] = 10'b0001000000;
assign label_6[420] = 10'b0001000000;
assign label_6[421] = 10'b0001000000;
assign label_6[422] = 10'b0000000100;
assign label_6[423] = 10'b0000000100;
assign label_6[424] = 10'b0000010000;
assign label_6[425] = 10'b0000010000;
assign label_6[426] = 10'b0000010000;
assign label_6[427] = 10'b0000010000;
assign label_6[428] = 10'b0001000000;
assign label_6[429] = 10'b0001000000;
assign label_6[430] = 10'b0001000000;
assign label_6[431] = 10'b0001000000;
assign label_6[432] = 10'b0100000000;
assign label_6[433] = 10'b0100000000;
assign label_6[434] = 10'b0100000000;
assign label_6[435] = 10'b0100000000;
assign label_6[436] = 10'b0100000000;
assign label_6[437] = 10'b0100000000;
assign label_6[438] = 10'b0100000000;
assign label_6[439] = 10'b0100000000;
assign label_6[440] = 10'b0000000100;
assign label_6[441] = 10'b0000000100;
assign label_6[442] = 10'b0000000100;
assign label_6[443] = 10'b0000000100;
assign label_6[444] = 10'b0000000100;
assign label_6[445] = 10'b0000000100;
assign label_6[446] = 10'b0000000100;
assign label_6[447] = 10'b0000000100;
assign label_6[448] = 10'b0010000000;
assign label_6[449] = 10'b0000001000;
assign label_6[450] = 10'b0000000100;
assign label_6[451] = 10'b0000000100;
assign label_6[452] = 10'b0100000000;
assign label_6[453] = 10'b0100000000;
assign label_6[454] = 10'b0000001000;
assign label_6[455] = 10'b0100000000;
assign label_6[456] = 10'b0000001000;
assign label_6[457] = 10'b0000000100;
assign label_6[458] = 10'b0010000000;
assign label_6[459] = 10'b0000000100;
assign label_6[460] = 10'b1000000000;
assign label_6[461] = 10'b1000000000;
assign label_6[462] = 10'b0010000000;
assign label_6[463] = 10'b1000000000;
assign label_6[464] = 10'b0000010000;
assign label_6[465] = 10'b1000000000;
assign label_6[466] = 10'b0000010000;
assign label_6[467] = 10'b0100000000;
assign label_6[468] = 10'b0000100000;
assign label_6[469] = 10'b0000100000;
assign label_6[470] = 10'b0000010000;
assign label_6[471] = 10'b0100000000;
assign label_6[472] = 10'b1000000000;
assign label_6[473] = 10'b0000000001;
assign label_6[474] = 10'b1000000000;
assign label_6[475] = 10'b0100000000;
assign label_6[476] = 10'b0000100000;
assign label_6[477] = 10'b0100000000;
assign label_6[478] = 10'b0100000000;
assign label_6[479] = 10'b0100000000;
assign label_6[480] = 10'b0000010000;
assign label_6[481] = 10'b1000000000;
assign label_6[482] = 10'b0000100000;
assign label_6[483] = 10'b1000000000;
assign label_6[484] = 10'b0000010000;
assign label_6[485] = 10'b1000000000;
assign label_6[486] = 10'b1000000000;
assign label_6[487] = 10'b1000000000;
assign label_6[488] = 10'b0000010000;
assign label_6[489] = 10'b1000000000;
assign label_6[490] = 10'b0000010000;
assign label_6[491] = 10'b1000000000;
assign label_6[492] = 10'b0000001000;
assign label_6[493] = 10'b0000100000;
assign label_6[494] = 10'b0000010000;
assign label_6[495] = 10'b0010000000;
assign label_6[496] = 10'b0000100000;
assign label_6[497] = 10'b0000100000;
assign label_6[498] = 10'b0000001000;
assign label_6[499] = 10'b0000001000;
assign label_6[500] = 10'b1000000000;
assign label_6[501] = 10'b0000100000;
assign label_6[502] = 10'b0000100000;
assign label_6[503] = 10'b1000000000;
assign label_6[504] = 10'b0000000001;
assign label_6[505] = 10'b0100000000;
assign label_6[506] = 10'b0100000000;
assign label_6[507] = 10'b0100000000;
assign label_6[508] = 10'b0001000000;
assign label_6[509] = 10'b0000000001;
assign label_6[510] = 10'b0001000000;
assign label_6[511] = 10'b0100000000;
assign label_6[512] = 10'b0000000001;
assign label_6[513] = 10'b0000000100;
assign label_6[514] = 10'b0000001000;
assign label_6[515] = 10'b0001000000;
assign label_6[516] = 10'b0000000100;
assign label_6[517] = 10'b0000000100;
assign label_6[518] = 10'b0000001000;
assign label_6[519] = 10'b0001000000;
assign label_6[520] = 10'b0000000001;
assign label_6[521] = 10'b0010000000;
assign label_6[522] = 10'b1000000000;
assign label_6[523] = 10'b0000001000;
assign label_6[524] = 10'b0000000001;
assign label_6[525] = 10'b0000010000;
assign label_6[526] = 10'b0000000001;
assign label_6[527] = 10'b1000000000;
assign label_6[528] = 10'b0000000010;
assign label_6[529] = 10'b0100000000;
assign label_6[530] = 10'b0100000000;
assign label_6[531] = 10'b0100000000;
assign label_6[532] = 10'b0000000100;
assign label_6[533] = 10'b0000000100;
assign label_6[534] = 10'b0000001000;
assign label_6[535] = 10'b0000001000;
assign label_6[536] = 10'b0000001000;
assign label_6[537] = 10'b0000001000;
assign label_6[538] = 10'b0100000000;
assign label_6[539] = 10'b0000000001;
assign label_6[540] = 10'b0000000010;
assign label_6[541] = 10'b0010000000;
assign label_6[542] = 10'b0000000010;
assign label_6[543] = 10'b0010000000;
assign label_6[544] = 10'b0000100000;
assign label_6[545] = 10'b0000000100;
assign label_6[546] = 10'b0000000100;
assign label_6[547] = 10'b0000000100;
assign label_6[548] = 10'b0000000100;
assign label_6[549] = 10'b0001000000;
assign label_6[550] = 10'b0000000100;
assign label_6[551] = 10'b0000000100;
assign label_6[552] = 10'b0000000100;
assign label_6[553] = 10'b0000010000;
assign label_6[554] = 10'b0001000000;
assign label_6[555] = 10'b0000010000;
assign label_6[556] = 10'b0001000000;
assign label_6[557] = 10'b0000000001;
assign label_6[558] = 10'b0000010000;
assign label_6[559] = 10'b0001000000;
assign label_6[560] = 10'b0000000100;
assign label_6[561] = 10'b0000000100;
assign label_6[562] = 10'b0100000000;
assign label_6[563] = 10'b0000100000;
assign label_6[564] = 10'b1000000000;
assign label_6[565] = 10'b0000000001;
assign label_6[566] = 10'b0010000000;
assign label_6[567] = 10'b0000000100;
assign label_6[568] = 10'b0000000100;
assign label_6[569] = 10'b0000001000;
assign label_6[570] = 10'b0000000100;
assign label_6[571] = 10'b0010000000;
assign label_6[572] = 10'b0010000000;
assign label_6[573] = 10'b0000000100;
assign label_6[574] = 10'b0000001000;
assign label_6[575] = 10'b0100000000;
assign label_6[576] = 10'b0000100000;
assign label_6[577] = 10'b0000000100;
assign label_6[578] = 10'b0000000001;
assign label_6[579] = 10'b0000000001;
assign label_6[580] = 10'b0100000000;
assign label_6[581] = 10'b0000100000;
assign label_6[582] = 10'b0100000000;
assign label_6[583] = 10'b0001000000;
assign label_6[584] = 10'b0000000001;
assign label_6[585] = 10'b0000100000;
assign label_6[586] = 10'b0000000001;
assign label_6[587] = 10'b0000001000;
assign label_6[588] = 10'b0001000000;
assign label_6[589] = 10'b0000010000;
assign label_6[590] = 10'b0000000100;
assign label_6[591] = 10'b0100000000;
assign label_6[592] = 10'b0001000000;
assign label_6[593] = 10'b0000100000;
assign label_6[594] = 10'b0000001000;
assign label_6[595] = 10'b0000000001;
assign label_6[596] = 10'b0001000000;
assign label_6[597] = 10'b0000000001;
assign label_6[598] = 10'b0000001000;
assign label_6[599] = 10'b0000000001;
assign label_6[600] = 10'b0001000000;
assign label_6[601] = 10'b0000000100;
assign label_6[602] = 10'b0000100000;
assign label_6[603] = 10'b0001000000;
assign label_6[604] = 10'b0000010000;
assign label_6[605] = 10'b0000100000;
assign label_6[606] = 10'b0000000100;
assign label_6[607] = 10'b0001000000;
assign label_6[608] = 10'b0100000000;
assign label_6[609] = 10'b0000100000;
assign label_6[610] = 10'b0000000001;
assign label_6[611] = 10'b0000001000;
assign label_6[612] = 10'b0000001000;
assign label_6[613] = 10'b0000001000;
assign label_6[614] = 10'b0000100000;
assign label_6[615] = 10'b0100000000;
assign label_6[616] = 10'b0000100000;
assign label_6[617] = 10'b0100000000;
assign label_6[618] = 10'b0000000001;
assign label_6[619] = 10'b0100000000;
assign label_6[620] = 10'b0100000000;
assign label_6[621] = 10'b0000001000;
assign label_6[622] = 10'b0000000001;
assign label_6[623] = 10'b0100000000;
assign label_6[624] = 10'b0000100000;
assign label_6[625] = 10'b0000001000;
assign label_6[626] = 10'b0000000001;
assign label_6[627] = 10'b0000000001;
assign label_6[628] = 10'b0000100000;
assign label_6[629] = 10'b0100000000;
assign label_6[630] = 10'b0000000001;
assign label_6[631] = 10'b0000010000;
assign label_6[632] = 10'b0000100000;
assign label_6[633] = 10'b0100000000;
assign label_6[634] = 10'b0000100000;
assign label_6[635] = 10'b0000000001;
assign label_6[636] = 10'b0000100000;
assign label_6[637] = 10'b0000000001;
assign label_6[638] = 10'b0000000001;
assign label_6[639] = 10'b0100000000;
assign label_6[640] = 10'b0000000100;
assign label_6[641] = 10'b0000001000;
assign label_6[642] = 10'b0000001000;
assign label_6[643] = 10'b0000000100;
assign label_6[644] = 10'b0000001000;
assign label_6[645] = 10'b0000000100;
assign label_6[646] = 10'b0000000100;
assign label_6[647] = 10'b0000000100;
assign label_6[648] = 10'b0000000100;
assign label_6[649] = 10'b0000000100;
assign label_6[650] = 10'b0100000000;
assign label_6[651] = 10'b0100000000;
assign label_6[652] = 10'b0000000100;
assign label_6[653] = 10'b0000000100;
assign label_6[654] = 10'b0000000100;
assign label_6[655] = 10'b0000000100;
assign label_6[656] = 10'b0000000100;
assign label_6[657] = 10'b0000010000;
assign label_6[658] = 10'b0000000100;
assign label_6[659] = 10'b0000000100;
assign label_6[660] = 10'b0000001000;
assign label_6[661] = 10'b0001000000;
assign label_6[662] = 10'b0000000100;
assign label_6[663] = 10'b0000000100;
assign label_6[664] = 10'b0000001000;
assign label_6[665] = 10'b0000001000;
assign label_6[666] = 10'b0000001000;
assign label_6[667] = 10'b0000001000;
assign label_6[668] = 10'b0000001000;
assign label_6[669] = 10'b0000001000;
assign label_6[670] = 10'b0000001000;
assign label_6[671] = 10'b0000001000;
assign label_6[672] = 10'b1000000000;
assign label_6[673] = 10'b1000000000;
assign label_6[674] = 10'b0000000001;
assign label_6[675] = 10'b0100000000;
assign label_6[676] = 10'b0100000000;
assign label_6[677] = 10'b0100000000;
assign label_6[678] = 10'b0100000000;
assign label_6[679] = 10'b0100000000;
assign label_6[680] = 10'b0100000000;
assign label_6[681] = 10'b0100000000;
assign label_6[682] = 10'b0000000100;
assign label_6[683] = 10'b0000000100;
assign label_6[684] = 10'b0100000000;
assign label_6[685] = 10'b0100000000;
assign label_6[686] = 10'b1000000000;
assign label_6[687] = 10'b1000000000;
assign label_6[688] = 10'b0000000100;
assign label_6[689] = 10'b0000000100;
assign label_6[690] = 10'b0000000100;
assign label_6[691] = 10'b0000000100;
assign label_6[692] = 10'b0001000000;
assign label_6[693] = 10'b0001000000;
assign label_6[694] = 10'b0001000000;
assign label_6[695] = 10'b0001000000;
assign label_6[696] = 10'b0000000001;
assign label_6[697] = 10'b0000000001;
assign label_6[698] = 10'b0001000000;
assign label_6[699] = 10'b0001000000;
assign label_6[700] = 10'b1000000000;
assign label_6[701] = 10'b1000000000;
assign label_6[702] = 10'b1000000000;
assign label_6[703] = 10'b0001000000;
assign label_6[704] = 10'b0000100000;
assign label_6[705] = 10'b0000000001;
assign label_6[706] = 10'b0000000100;
assign label_6[707] = 10'b0000001000;
assign label_6[708] = 10'b0000000001;
assign label_6[709] = 10'b0000000100;
assign label_6[710] = 10'b0000001000;
assign label_6[711] = 10'b0000001000;
assign label_6[712] = 10'b0000001000;
assign label_6[713] = 10'b0000000100;
assign label_6[714] = 10'b0000100000;
assign label_6[715] = 10'b0000100000;
assign label_6[716] = 10'b0000001000;
assign label_6[717] = 10'b0000000100;
assign label_6[718] = 10'b0000000100;
assign label_6[719] = 10'b0000000100;
assign label_6[720] = 10'b0000001000;
assign label_6[721] = 10'b0000001000;
assign label_6[722] = 10'b0000001000;
assign label_6[723] = 10'b0000000100;
assign label_6[724] = 10'b0000001000;
assign label_6[725] = 10'b0000001000;
assign label_6[726] = 10'b0000000001;
assign label_6[727] = 10'b0000001000;
assign label_6[728] = 10'b0000100000;
assign label_6[729] = 10'b0100000000;
assign label_6[730] = 10'b0000100000;
assign label_6[731] = 10'b0000001000;
assign label_6[732] = 10'b0000100000;
assign label_6[733] = 10'b0000001000;
assign label_6[734] = 10'b0000001000;
assign label_6[735] = 10'b0000001000;
assign label_6[736] = 10'b0000000100;
assign label_6[737] = 10'b0100000000;
assign label_6[738] = 10'b0000000100;
assign label_6[739] = 10'b0000001000;
assign label_6[740] = 10'b0000000100;
assign label_6[741] = 10'b0000001000;
assign label_6[742] = 10'b0000000100;
assign label_6[743] = 10'b0100000000;
assign label_6[744] = 10'b0000001000;
assign label_6[745] = 10'b0100000000;
assign label_6[746] = 10'b0000001000;
assign label_6[747] = 10'b0000001000;
assign label_6[748] = 10'b0000000100;
assign label_6[749] = 10'b0000000100;
assign label_6[750] = 10'b0100000000;
assign label_6[751] = 10'b0000001000;
assign label_6[752] = 10'b0000000100;
assign label_6[753] = 10'b0000000100;
assign label_6[754] = 10'b0000000100;
assign label_6[755] = 10'b0100000000;
assign label_6[756] = 10'b0001000000;
assign label_6[757] = 10'b0000100000;
assign label_6[758] = 10'b0000100000;
assign label_6[759] = 10'b0000000001;
assign label_6[760] = 10'b0000001000;
assign label_6[761] = 10'b0000001000;
assign label_6[762] = 10'b0000100000;
assign label_6[763] = 10'b0100000000;
assign label_6[764] = 10'b0100000000;
assign label_6[765] = 10'b0000000100;
assign label_6[766] = 10'b0100000000;
assign label_6[767] = 10'b0000000100;
assign label_6[768] = 10'b0000000001;
assign label_6[769] = 10'b0000010000;
assign label_6[770] = 10'b0000100000;
assign label_6[771] = 10'b0000100000;
assign label_6[772] = 10'b0000100000;
assign label_6[773] = 10'b0000100000;
assign label_6[774] = 10'b0001000000;
assign label_6[775] = 10'b0001000000;
assign label_6[776] = 10'b0000100000;
assign label_6[777] = 10'b1000000000;
assign label_6[778] = 10'b0000010000;
assign label_6[779] = 10'b0001000000;
assign label_6[780] = 10'b0001000000;
assign label_6[781] = 10'b0001000000;
assign label_6[782] = 10'b0000000001;
assign label_6[783] = 10'b0000010000;
assign label_6[784] = 10'b1000000000;
assign label_6[785] = 10'b0001000000;
assign label_6[786] = 10'b0000010000;
assign label_6[787] = 10'b1000000000;
assign label_6[788] = 10'b0001000000;
assign label_6[789] = 10'b0001000000;
assign label_6[790] = 10'b0000010000;
assign label_6[791] = 10'b0001000000;
assign label_6[792] = 10'b0000010000;
assign label_6[793] = 10'b0000010000;
assign label_6[794] = 10'b0000000100;
assign label_6[795] = 10'b0000000001;
assign label_6[796] = 10'b1000000000;
assign label_6[797] = 10'b0000000100;
assign label_6[798] = 10'b0000000001;
assign label_6[799] = 10'b0100000000;
assign label_6[800] = 10'b0000100000;
assign label_6[801] = 10'b0000010000;
assign label_6[802] = 10'b0000000100;
assign label_6[803] = 10'b0000000100;
assign label_6[804] = 10'b0000000100;
assign label_6[805] = 10'b0010000000;
assign label_6[806] = 10'b0000010000;
assign label_6[807] = 10'b1000000000;
assign label_6[808] = 10'b0000000001;
assign label_6[809] = 10'b0000000001;
assign label_6[810] = 10'b0000000001;
assign label_6[811] = 10'b0000000001;
assign label_6[812] = 10'b0000100000;
assign label_6[813] = 10'b0000100000;
assign label_6[814] = 10'b0000100000;
assign label_6[815] = 10'b0000100000;
assign label_6[816] = 10'b0000000001;
assign label_6[817] = 10'b1000000000;
assign label_6[818] = 10'b0010000000;
assign label_6[819] = 10'b0001000000;
assign label_6[820] = 10'b0000000001;
assign label_6[821] = 10'b0000000001;
assign label_6[822] = 10'b0001000000;
assign label_6[823] = 10'b0001000000;
assign label_6[824] = 10'b0000000001;
assign label_6[825] = 10'b0000010000;
assign label_6[826] = 10'b0000000100;
assign label_6[827] = 10'b1000000000;
assign label_6[828] = 10'b0000000001;
assign label_6[829] = 10'b0001000000;
assign label_6[830] = 10'b0000000001;
assign label_6[831] = 10'b0000000001;
assign label_6[832] = 10'b0000100000;
assign label_6[833] = 10'b0000000100;
assign label_6[834] = 10'b0000000001;
assign label_6[835] = 10'b1000000000;
assign label_6[836] = 10'b0000000001;
assign label_6[837] = 10'b0000100000;
assign label_6[838] = 10'b0001000000;
assign label_6[839] = 10'b0100000000;
assign label_6[840] = 10'b0000100000;
assign label_6[841] = 10'b0000100000;
assign label_6[842] = 10'b0000100000;
assign label_6[843] = 10'b0000100000;
assign label_6[844] = 10'b0000000001;
assign label_6[845] = 10'b0000000001;
assign label_6[846] = 10'b0000100000;
assign label_6[847] = 10'b0000000001;
assign label_6[848] = 10'b0000100000;
assign label_6[849] = 10'b0000001000;
assign label_6[850] = 10'b0000001000;
assign label_6[851] = 10'b0000000100;
assign label_6[852] = 10'b0000100000;
assign label_6[853] = 10'b0000001000;
assign label_6[854] = 10'b0000000001;
assign label_6[855] = 10'b0000100000;
assign label_6[856] = 10'b0000000100;
assign label_6[857] = 10'b0000000100;
assign label_6[858] = 10'b0000000001;
assign label_6[859] = 10'b0000100000;
assign label_6[860] = 10'b0000000001;
assign label_6[861] = 10'b0000000001;
assign label_6[862] = 10'b0100000000;
assign label_6[863] = 10'b0000000001;
assign label_6[864] = 10'b0000100000;
assign label_6[865] = 10'b0000001000;
assign label_6[866] = 10'b0000000001;
assign label_6[867] = 10'b0000100000;
assign label_6[868] = 10'b0000000001;
assign label_6[869] = 10'b0000000001;
assign label_6[870] = 10'b0000100000;
assign label_6[871] = 10'b0000000001;
assign label_6[872] = 10'b0001000000;
assign label_6[873] = 10'b0000000001;
assign label_6[874] = 10'b0000000001;
assign label_6[875] = 10'b0000000100;
assign label_6[876] = 10'b0000000100;
assign label_6[877] = 10'b0001000000;
assign label_6[878] = 10'b1000000000;
assign label_6[879] = 10'b1000000000;
assign label_6[880] = 10'b0100000000;
assign label_6[881] = 10'b0100000000;
assign label_6[882] = 10'b0100000000;
assign label_6[883] = 10'b0100000000;
assign label_6[884] = 10'b0000100000;
assign label_6[885] = 10'b0000010000;
assign label_6[886] = 10'b0001000000;
assign label_6[887] = 10'b0000000100;
assign label_6[888] = 10'b0000000001;
assign label_6[889] = 10'b0001000000;
assign label_6[890] = 10'b0001000000;
assign label_6[891] = 10'b0000000100;
assign label_6[892] = 10'b0000000001;
assign label_6[893] = 10'b0100000000;
assign label_6[894] = 10'b0000000001;
assign label_6[895] = 10'b0000000001;
assign label_6[896] = 10'b0000100000;
assign label_6[897] = 10'b0001000000;
assign label_6[898] = 10'b0000001000;
assign label_6[899] = 10'b0000100000;
assign label_6[900] = 10'b0000000100;
assign label_6[901] = 10'b0000000100;
assign label_6[902] = 10'b0001000000;
assign label_6[903] = 10'b0000000100;
assign label_6[904] = 10'b0001000000;
assign label_6[905] = 10'b0001000000;
assign label_6[906] = 10'b0001000000;
assign label_6[907] = 10'b0001000000;
assign label_6[908] = 10'b0000000001;
assign label_6[909] = 10'b0000000001;
assign label_6[910] = 10'b0000000001;
assign label_6[911] = 10'b0000000001;
assign label_6[912] = 10'b0000001000;
assign label_6[913] = 10'b0000100000;
assign label_6[914] = 10'b0000100000;
assign label_6[915] = 10'b0000001000;
assign label_6[916] = 10'b0000100000;
assign label_6[917] = 10'b0000100000;
assign label_6[918] = 10'b0000000001;
assign label_6[919] = 10'b0000001000;
assign label_6[920] = 10'b0000010000;
assign label_6[921] = 10'b0000100000;
assign label_6[922] = 10'b0100000000;
assign label_6[923] = 10'b0000001000;
assign label_6[924] = 10'b0000001000;
assign label_6[925] = 10'b0000100000;
assign label_6[926] = 10'b0000001000;
assign label_6[927] = 10'b0000000100;
assign label_6[928] = 10'b0000100000;
assign label_6[929] = 10'b0000100000;
assign label_6[930] = 10'b0100000000;
assign label_6[931] = 10'b0000000100;
assign label_6[932] = 10'b1000000000;
assign label_6[933] = 10'b0100000000;
assign label_6[934] = 10'b0000001000;
assign label_6[935] = 10'b0000010000;
assign label_6[936] = 10'b0000001000;
assign label_6[937] = 10'b0000100000;
assign label_6[938] = 10'b0000001000;
assign label_6[939] = 10'b0000001000;
assign label_6[940] = 10'b0000000100;
assign label_6[941] = 10'b0000010000;
assign label_6[942] = 10'b0001000000;
assign label_6[943] = 10'b0100000000;
assign label_6[944] = 10'b0100000000;
assign label_6[945] = 10'b0001000000;
assign label_6[946] = 10'b0000000100;
assign label_6[947] = 10'b0000010000;
assign label_6[948] = 10'b0100000000;
assign label_6[949] = 10'b0000000100;
assign label_6[950] = 10'b0000000100;
assign label_6[951] = 10'b0001000000;
assign label_6[952] = 10'b0000000001;
assign label_6[953] = 10'b0000100000;
assign label_6[954] = 10'b0000000001;
assign label_6[955] = 10'b0001000000;
assign label_6[956] = 10'b0001000000;
assign label_6[957] = 10'b0001000000;
assign label_6[958] = 10'b0001000000;
assign label_6[959] = 10'b0001000000;
assign label_6[960] = 10'b0000001000;
assign label_6[961] = 10'b0100000000;
assign label_6[962] = 10'b0001000000;
assign label_6[963] = 10'b0000100000;
assign label_6[964] = 10'b0000000100;
assign label_6[965] = 10'b0001000000;
assign label_6[966] = 10'b0000001000;
assign label_6[967] = 10'b0000000100;
assign label_6[968] = 10'b0000000100;
assign label_6[969] = 10'b0000000100;
assign label_6[970] = 10'b0000000001;
assign label_6[971] = 10'b0000100000;
assign label_6[972] = 10'b0000100000;
assign label_6[973] = 10'b0100000000;
assign label_6[974] = 10'b0000100000;
assign label_6[975] = 10'b0100000000;
assign label_6[976] = 10'b0000000100;
assign label_6[977] = 10'b0000001000;
assign label_6[978] = 10'b0001000000;
assign label_6[979] = 10'b0001000000;
assign label_6[980] = 10'b0000100000;
assign label_6[981] = 10'b0000100000;
assign label_6[982] = 10'b0000100000;
assign label_6[983] = 10'b0000100000;
assign label_6[984] = 10'b0001000000;
assign label_6[985] = 10'b0001000000;
assign label_6[986] = 10'b0000000100;
assign label_6[987] = 10'b0000000100;
assign label_6[988] = 10'b0001000000;
assign label_6[989] = 10'b0001000000;
assign label_6[990] = 10'b0000100000;
assign label_6[991] = 10'b0001000000;
assign label_6[992] = 10'b0000010000;
assign label_6[993] = 10'b0100000000;
assign label_6[994] = 10'b0001000000;
assign label_6[995] = 10'b0100000000;
assign label_6[996] = 10'b1000000000;
assign label_6[997] = 10'b0100000000;
assign label_6[998] = 10'b0000100000;
assign label_6[999] = 10'b0100000000;
assign label_6[1000] = 10'b0000100000;
assign label_6[1001] = 10'b0000000100;
assign label_6[1002] = 10'b0000100000;
assign label_6[1003] = 10'b0100000000;
assign label_6[1004] = 10'b0001000000;
assign label_6[1005] = 10'b0000010000;
assign label_6[1006] = 10'b0000010000;
assign label_6[1007] = 10'b0000000001;
assign label_6[1008] = 10'b0000001000;
assign label_6[1009] = 10'b0000000100;
assign label_6[1010] = 10'b0100000000;
assign label_6[1011] = 10'b0100000000;
assign label_6[1012] = 10'b0100000000;
assign label_6[1013] = 10'b0100000000;
assign label_6[1014] = 10'b0000000100;
assign label_6[1015] = 10'b0100000000;
assign label_6[1016] = 10'b0000000100;
assign label_6[1017] = 10'b0000000001;
assign label_6[1018] = 10'b0100000000;
assign label_6[1019] = 10'b0000000001;
assign label_6[1020] = 10'b0000010000;
assign label_6[1021] = 10'b0000010000;
assign label_6[1022] = 10'b0100000000;
assign label_6[1023] = 10'b0100000000;
assign label_7[0] = 10'b0010000000;
assign label_7[1] = 10'b0000000001;
assign label_7[2] = 10'b1000000000;
assign label_7[3] = 10'b0010000000;
assign label_7[4] = 10'b0000010000;
assign label_7[5] = 10'b0000010000;
assign label_7[6] = 10'b0000100000;
assign label_7[7] = 10'b1000000000;
assign label_7[8] = 10'b0010000000;
assign label_7[9] = 10'b0000000001;
assign label_7[10] = 10'b0001000000;
assign label_7[11] = 10'b0001000000;
assign label_7[12] = 10'b0000000001;
assign label_7[13] = 10'b0000000001;
assign label_7[14] = 10'b0000000001;
assign label_7[15] = 10'b0000000001;
assign label_7[16] = 10'b0010000000;
assign label_7[17] = 10'b1000000000;
assign label_7[18] = 10'b0000001000;
assign label_7[19] = 10'b0000010000;
assign label_7[20] = 10'b0000010000;
assign label_7[21] = 10'b1000000000;
assign label_7[22] = 10'b0000010000;
assign label_7[23] = 10'b1000000000;
assign label_7[24] = 10'b0010000000;
assign label_7[25] = 10'b1000000000;
assign label_7[26] = 10'b0000001000;
assign label_7[27] = 10'b0000000010;
assign label_7[28] = 10'b1000000000;
assign label_7[29] = 10'b0000001000;
assign label_7[30] = 10'b0000000010;
assign label_7[31] = 10'b1000000000;
assign label_7[32] = 10'b0010000000;
assign label_7[33] = 10'b0000100000;
assign label_7[34] = 10'b0000010000;
assign label_7[35] = 10'b0010000000;
assign label_7[36] = 10'b0000010000;
assign label_7[37] = 10'b1000000000;
assign label_7[38] = 10'b1000000000;
assign label_7[39] = 10'b1000000000;
assign label_7[40] = 10'b0000100000;
assign label_7[41] = 10'b0001000000;
assign label_7[42] = 10'b0001000000;
assign label_7[43] = 10'b0000010000;
assign label_7[44] = 10'b0000001000;
assign label_7[45] = 10'b0000001000;
assign label_7[46] = 10'b0000001000;
assign label_7[47] = 10'b0000001000;
assign label_7[48] = 10'b0000100000;
assign label_7[49] = 10'b0000100000;
assign label_7[50] = 10'b0000001000;
assign label_7[51] = 10'b0000100000;
assign label_7[52] = 10'b0000001000;
assign label_7[53] = 10'b0000100000;
assign label_7[54] = 10'b0000001000;
assign label_7[55] = 10'b0000100000;
assign label_7[56] = 10'b1000000000;
assign label_7[57] = 10'b0000100000;
assign label_7[58] = 10'b0000000001;
assign label_7[59] = 10'b0000000001;
assign label_7[60] = 10'b0000100000;
assign label_7[61] = 10'b0000100000;
assign label_7[62] = 10'b0000001000;
assign label_7[63] = 10'b0000001000;
assign label_7[64] = 10'b0001000000;
assign label_7[65] = 10'b1000000000;
assign label_7[66] = 10'b0000100000;
assign label_7[67] = 10'b0000010000;
assign label_7[68] = 10'b0001000000;
assign label_7[69] = 10'b0001000000;
assign label_7[70] = 10'b0000010000;
assign label_7[71] = 10'b0100000000;
assign label_7[72] = 10'b1000000000;
assign label_7[73] = 10'b0000000001;
assign label_7[74] = 10'b0001000000;
assign label_7[75] = 10'b0000000100;
assign label_7[76] = 10'b0001000000;
assign label_7[77] = 10'b0001000000;
assign label_7[78] = 10'b0000000001;
assign label_7[79] = 10'b0001000000;
assign label_7[80] = 10'b0000010000;
assign label_7[81] = 10'b1000000000;
assign label_7[82] = 10'b1000000000;
assign label_7[83] = 10'b0000000001;
assign label_7[84] = 10'b0000100000;
assign label_7[85] = 10'b0000010000;
assign label_7[86] = 10'b0000000001;
assign label_7[87] = 10'b0000010000;
assign label_7[88] = 10'b0001000000;
assign label_7[89] = 10'b0100000000;
assign label_7[90] = 10'b0100000000;
assign label_7[91] = 10'b0000100000;
assign label_7[92] = 10'b0000100000;
assign label_7[93] = 10'b0100000000;
assign label_7[94] = 10'b0000100000;
assign label_7[95] = 10'b0000000001;
assign label_7[96] = 10'b0001000000;
assign label_7[97] = 10'b0000000001;
assign label_7[98] = 10'b0001000000;
assign label_7[99] = 10'b0001000000;
assign label_7[100] = 10'b0000000100;
assign label_7[101] = 10'b0000000100;
assign label_7[102] = 10'b0000000010;
assign label_7[103] = 10'b0001000000;
assign label_7[104] = 10'b0000000100;
assign label_7[105] = 10'b0000000100;
assign label_7[106] = 10'b0000100000;
assign label_7[107] = 10'b0000100000;
assign label_7[108] = 10'b0000000001;
assign label_7[109] = 10'b0001000000;
assign label_7[110] = 10'b0001000000;
assign label_7[111] = 10'b0001000000;
assign label_7[112] = 10'b0000000100;
assign label_7[113] = 10'b0000000100;
assign label_7[114] = 10'b0000000100;
assign label_7[115] = 10'b0000000100;
assign label_7[116] = 10'b0000000100;
assign label_7[117] = 10'b0000000100;
assign label_7[118] = 10'b0000000100;
assign label_7[119] = 10'b0000000100;
assign label_7[120] = 10'b0000000100;
assign label_7[121] = 10'b0000000100;
assign label_7[122] = 10'b0000000100;
assign label_7[123] = 10'b0000000100;
assign label_7[124] = 10'b0000000100;
assign label_7[125] = 10'b0000000100;
assign label_7[126] = 10'b0000000100;
assign label_7[127] = 10'b0000000100;
assign label_7[128] = 10'b0000000100;
assign label_7[129] = 10'b0000001000;
assign label_7[130] = 10'b0001000000;
assign label_7[131] = 10'b0000001000;
assign label_7[132] = 10'b0000010000;
assign label_7[133] = 10'b0000000010;
assign label_7[134] = 10'b0000001000;
assign label_7[135] = 10'b0000010000;
assign label_7[136] = 10'b0000001000;
assign label_7[137] = 10'b0000000100;
assign label_7[138] = 10'b0000100000;
assign label_7[139] = 10'b0000001000;
assign label_7[140] = 10'b0000000100;
assign label_7[141] = 10'b0100000000;
assign label_7[142] = 10'b0000000100;
assign label_7[143] = 10'b0001000000;
assign label_7[144] = 10'b0000001000;
assign label_7[145] = 10'b0000000100;
assign label_7[146] = 10'b0000001000;
assign label_7[147] = 10'b0000001000;
assign label_7[148] = 10'b0000100000;
assign label_7[149] = 10'b0000001000;
assign label_7[150] = 10'b0000100000;
assign label_7[151] = 10'b0000001000;
assign label_7[152] = 10'b0100000000;
assign label_7[153] = 10'b0100000000;
assign label_7[154] = 10'b0000000001;
assign label_7[155] = 10'b0000100000;
assign label_7[156] = 10'b0000001000;
assign label_7[157] = 10'b0000100000;
assign label_7[158] = 10'b0000000100;
assign label_7[159] = 10'b0000001000;
assign label_7[160] = 10'b0000100000;
assign label_7[161] = 10'b0001000000;
assign label_7[162] = 10'b0100000000;
assign label_7[163] = 10'b0000000001;
assign label_7[164] = 10'b0001000000;
assign label_7[165] = 10'b0000100000;
assign label_7[166] = 10'b0000000001;
assign label_7[167] = 10'b0100000000;
assign label_7[168] = 10'b0000100000;
assign label_7[169] = 10'b0100000000;
assign label_7[170] = 10'b0000000100;
assign label_7[171] = 10'b0000001000;
assign label_7[172] = 10'b0100000000;
assign label_7[173] = 10'b0000000100;
assign label_7[174] = 10'b0001000000;
assign label_7[175] = 10'b0100000000;
assign label_7[176] = 10'b0000000010;
assign label_7[177] = 10'b0000001000;
assign label_7[178] = 10'b0000001000;
assign label_7[179] = 10'b0000001000;
assign label_7[180] = 10'b0100000000;
assign label_7[181] = 10'b0000000010;
assign label_7[182] = 10'b0000001000;
assign label_7[183] = 10'b0000100000;
assign label_7[184] = 10'b0000000100;
assign label_7[185] = 10'b0000100000;
assign label_7[186] = 10'b0100000000;
assign label_7[187] = 10'b0100000000;
assign label_7[188] = 10'b0000000001;
assign label_7[189] = 10'b0100000000;
assign label_7[190] = 10'b0000000001;
assign label_7[191] = 10'b0000001000;
assign label_7[192] = 10'b0001000000;
assign label_7[193] = 10'b0000000100;
assign label_7[194] = 10'b0001000000;
assign label_7[195] = 10'b0000100000;
assign label_7[196] = 10'b0000000001;
assign label_7[197] = 10'b0000000001;
assign label_7[198] = 10'b0000000100;
assign label_7[199] = 10'b0000000100;
assign label_7[200] = 10'b0000000001;
assign label_7[201] = 10'b0000010000;
assign label_7[202] = 10'b0000000100;
assign label_7[203] = 10'b1000000000;
assign label_7[204] = 10'b0000010000;
assign label_7[205] = 10'b0000000001;
assign label_7[206] = 10'b0100000000;
assign label_7[207] = 10'b0000010000;
assign label_7[208] = 10'b0000000001;
assign label_7[209] = 10'b0000000001;
assign label_7[210] = 10'b0000100000;
assign label_7[211] = 10'b0000100000;
assign label_7[212] = 10'b0000000001;
assign label_7[213] = 10'b0001000000;
assign label_7[214] = 10'b0000000001;
assign label_7[215] = 10'b0000010000;
assign label_7[216] = 10'b0000100000;
assign label_7[217] = 10'b0000100000;
assign label_7[218] = 10'b0000000001;
assign label_7[219] = 10'b0000001000;
assign label_7[220] = 10'b0000100000;
assign label_7[221] = 10'b0001000000;
assign label_7[222] = 10'b0000100000;
assign label_7[223] = 10'b0000000001;
assign label_7[224] = 10'b0000000100;
assign label_7[225] = 10'b0000100000;
assign label_7[226] = 10'b0100000000;
assign label_7[227] = 10'b0000001000;
assign label_7[228] = 10'b0000000100;
assign label_7[229] = 10'b0001000000;
assign label_7[230] = 10'b0001000000;
assign label_7[231] = 10'b0001000000;
assign label_7[232] = 10'b0000010000;
assign label_7[233] = 10'b0001000000;
assign label_7[234] = 10'b0000001000;
assign label_7[235] = 10'b0000000100;
assign label_7[236] = 10'b0000001000;
assign label_7[237] = 10'b0000001000;
assign label_7[238] = 10'b0000001000;
assign label_7[239] = 10'b0000000001;
assign label_7[240] = 10'b0000100000;
assign label_7[241] = 10'b0000000100;
assign label_7[242] = 10'b0000001000;
assign label_7[243] = 10'b0000100000;
assign label_7[244] = 10'b0000010000;
assign label_7[245] = 10'b1000000000;
assign label_7[246] = 10'b0000001000;
assign label_7[247] = 10'b0000000001;
assign label_7[248] = 10'b0000100000;
assign label_7[249] = 10'b0100000000;
assign label_7[250] = 10'b0001000000;
assign label_7[251] = 10'b0000000100;
assign label_7[252] = 10'b0000100000;
assign label_7[253] = 10'b0000000001;
assign label_7[254] = 10'b0100000000;
assign label_7[255] = 10'b0000000001;
assign label_7[256] = 10'b0000100000;
assign label_7[257] = 10'b0000001000;
assign label_7[258] = 10'b0000000100;
assign label_7[259] = 10'b0000001000;
assign label_7[260] = 10'b0000001000;
assign label_7[261] = 10'b0000000100;
assign label_7[262] = 10'b0000001000;
assign label_7[263] = 10'b0000001000;
assign label_7[264] = 10'b0000001000;
assign label_7[265] = 10'b0000001000;
assign label_7[266] = 10'b0000001000;
assign label_7[267] = 10'b0000000100;
assign label_7[268] = 10'b0000000100;
assign label_7[269] = 10'b0000000100;
assign label_7[270] = 10'b0000000100;
assign label_7[271] = 10'b0000001000;
assign label_7[272] = 10'b0000001000;
assign label_7[273] = 10'b0000100000;
assign label_7[274] = 10'b0000000001;
assign label_7[275] = 10'b0000000001;
assign label_7[276] = 10'b0000100000;
assign label_7[277] = 10'b0000000001;
assign label_7[278] = 10'b0100000000;
assign label_7[279] = 10'b0000001000;
assign label_7[280] = 10'b0000001000;
assign label_7[281] = 10'b0000100000;
assign label_7[282] = 10'b0000100000;
assign label_7[283] = 10'b0000001000;
assign label_7[284] = 10'b0000001000;
assign label_7[285] = 10'b0000100000;
assign label_7[286] = 10'b0100000000;
assign label_7[287] = 10'b0000000100;
assign label_7[288] = 10'b0000000100;
assign label_7[289] = 10'b0000100000;
assign label_7[290] = 10'b0000000100;
assign label_7[291] = 10'b0000000100;
assign label_7[292] = 10'b0000001000;
assign label_7[293] = 10'b0000100000;
assign label_7[294] = 10'b0100000000;
assign label_7[295] = 10'b0100000000;
assign label_7[296] = 10'b0000000100;
assign label_7[297] = 10'b0000000100;
assign label_7[298] = 10'b0001000000;
assign label_7[299] = 10'b0001000000;
assign label_7[300] = 10'b0000001000;
assign label_7[301] = 10'b0000100000;
assign label_7[302] = 10'b0000000100;
assign label_7[303] = 10'b0100000000;
assign label_7[304] = 10'b0000100000;
assign label_7[305] = 10'b0000100000;
assign label_7[306] = 10'b0001000000;
assign label_7[307] = 10'b0000000001;
assign label_7[308] = 10'b0001000000;
assign label_7[309] = 10'b0000000100;
assign label_7[310] = 10'b0000100000;
assign label_7[311] = 10'b0100000000;
assign label_7[312] = 10'b0000000001;
assign label_7[313] = 10'b0000000001;
assign label_7[314] = 10'b0000000001;
assign label_7[315] = 10'b0100000000;
assign label_7[316] = 10'b0000000100;
assign label_7[317] = 10'b0000000100;
assign label_7[318] = 10'b0000001000;
assign label_7[319] = 10'b0000001000;
assign label_7[320] = 10'b0000100000;
assign label_7[321] = 10'b0000000001;
assign label_7[322] = 10'b0000000100;
assign label_7[323] = 10'b0000000001;
assign label_7[324] = 10'b0000100000;
assign label_7[325] = 10'b0001000000;
assign label_7[326] = 10'b0000000001;
assign label_7[327] = 10'b0000000001;
assign label_7[328] = 10'b0000000001;
assign label_7[329] = 10'b0000000001;
assign label_7[330] = 10'b0000000001;
assign label_7[331] = 10'b0000100000;
assign label_7[332] = 10'b0001000000;
assign label_7[333] = 10'b0001000000;
assign label_7[334] = 10'b0001000000;
assign label_7[335] = 10'b0001000000;
assign label_7[336] = 10'b0000000001;
assign label_7[337] = 10'b0000010000;
assign label_7[338] = 10'b1000000000;
assign label_7[339] = 10'b0000000001;
assign label_7[340] = 10'b0000000001;
assign label_7[341] = 10'b0000000001;
assign label_7[342] = 10'b0010000000;
assign label_7[343] = 10'b0001000000;
assign label_7[344] = 10'b0000000001;
assign label_7[345] = 10'b0000000001;
assign label_7[346] = 10'b0000000100;
assign label_7[347] = 10'b0000000100;
assign label_7[348] = 10'b0000000001;
assign label_7[349] = 10'b0000000001;
assign label_7[350] = 10'b0001000000;
assign label_7[351] = 10'b0000000100;
assign label_7[352] = 10'b0000100000;
assign label_7[353] = 10'b0000100000;
assign label_7[354] = 10'b0000100000;
assign label_7[355] = 10'b0000001000;
assign label_7[356] = 10'b0000001000;
assign label_7[357] = 10'b0000100000;
assign label_7[358] = 10'b0000001000;
assign label_7[359] = 10'b0000000100;
assign label_7[360] = 10'b0000100000;
assign label_7[361] = 10'b0000001000;
assign label_7[362] = 10'b0000100000;
assign label_7[363] = 10'b0000000100;
assign label_7[364] = 10'b0000100000;
assign label_7[365] = 10'b0000000100;
assign label_7[366] = 10'b0000001000;
assign label_7[367] = 10'b0000001000;
assign label_7[368] = 10'b0000100000;
assign label_7[369] = 10'b0001000000;
assign label_7[370] = 10'b0001000000;
assign label_7[371] = 10'b0000100000;
assign label_7[372] = 10'b0000000100;
assign label_7[373] = 10'b0000000001;
assign label_7[374] = 10'b0000100000;
assign label_7[375] = 10'b0000100000;
assign label_7[376] = 10'b0000000001;
assign label_7[377] = 10'b0100000000;
assign label_7[378] = 10'b0000010000;
assign label_7[379] = 10'b0100000000;
assign label_7[380] = 10'b0000001000;
assign label_7[381] = 10'b0000000001;
assign label_7[382] = 10'b0000000100;
assign label_7[383] = 10'b0000000001;
assign label_7[384] = 10'b0000100000;
assign label_7[385] = 10'b0000001000;
assign label_7[386] = 10'b0000000001;
assign label_7[387] = 10'b0001000000;
assign label_7[388] = 10'b0000000001;
assign label_7[389] = 10'b0001000000;
assign label_7[390] = 10'b0001000000;
assign label_7[391] = 10'b0000000100;
assign label_7[392] = 10'b0001000000;
assign label_7[393] = 10'b0000010000;
assign label_7[394] = 10'b0000001000;
assign label_7[395] = 10'b0000100000;
assign label_7[396] = 10'b0000000001;
assign label_7[397] = 10'b0000000001;
assign label_7[398] = 10'b0001000000;
assign label_7[399] = 10'b0001000000;
assign label_7[400] = 10'b0000000001;
assign label_7[401] = 10'b0001000000;
assign label_7[402] = 10'b0000000100;
assign label_7[403] = 10'b0000001000;
assign label_7[404] = 10'b0000000001;
assign label_7[405] = 10'b0000000001;
assign label_7[406] = 10'b0100000000;
assign label_7[407] = 10'b0000000001;
assign label_7[408] = 10'b0000000100;
assign label_7[409] = 10'b0000000100;
assign label_7[410] = 10'b0000000100;
assign label_7[411] = 10'b0000000100;
assign label_7[412] = 10'b0000000100;
assign label_7[413] = 10'b0000000100;
assign label_7[414] = 10'b0000000100;
assign label_7[415] = 10'b0000000100;
assign label_7[416] = 10'b0000000001;
assign label_7[417] = 10'b0001000000;
assign label_7[418] = 10'b0000100000;
assign label_7[419] = 10'b0000001000;
assign label_7[420] = 10'b0000000100;
assign label_7[421] = 10'b0000001000;
assign label_7[422] = 10'b0000001000;
assign label_7[423] = 10'b0000100000;
assign label_7[424] = 10'b0100000000;
assign label_7[425] = 10'b0000100000;
assign label_7[426] = 10'b0000001000;
assign label_7[427] = 10'b0000001000;
assign label_7[428] = 10'b0000001000;
assign label_7[429] = 10'b0000000100;
assign label_7[430] = 10'b0000000100;
assign label_7[431] = 10'b0000000100;
assign label_7[432] = 10'b0000000001;
assign label_7[433] = 10'b0000001000;
assign label_7[434] = 10'b0000000100;
assign label_7[435] = 10'b0000010000;
assign label_7[436] = 10'b0000001000;
assign label_7[437] = 10'b0000001000;
assign label_7[438] = 10'b0000000001;
assign label_7[439] = 10'b0000000100;
assign label_7[440] = 10'b0000000001;
assign label_7[441] = 10'b0000001000;
assign label_7[442] = 10'b0000000100;
assign label_7[443] = 10'b0000001000;
assign label_7[444] = 10'b0000000001;
assign label_7[445] = 10'b0000000001;
assign label_7[446] = 10'b0000001000;
assign label_7[447] = 10'b0000001000;
assign label_7[448] = 10'b0000000001;
assign label_7[449] = 10'b0000000001;
assign label_7[450] = 10'b0000000001;
assign label_7[451] = 10'b0000010000;
assign label_7[452] = 10'b0001000000;
assign label_7[453] = 10'b0000010000;
assign label_7[454] = 10'b1000000000;
assign label_7[455] = 10'b0000000001;
assign label_7[456] = 10'b0001000000;
assign label_7[457] = 10'b0001000000;
assign label_7[458] = 10'b0001000000;
assign label_7[459] = 10'b0001000000;
assign label_7[460] = 10'b0000000001;
assign label_7[461] = 10'b0000000001;
assign label_7[462] = 10'b0000000001;
assign label_7[463] = 10'b0000000001;
assign label_7[464] = 10'b0001000000;
assign label_7[465] = 10'b0000000001;
assign label_7[466] = 10'b0000000001;
assign label_7[467] = 10'b0000010000;
assign label_7[468] = 10'b0001000000;
assign label_7[469] = 10'b0001000000;
assign label_7[470] = 10'b0001000000;
assign label_7[471] = 10'b0001000000;
assign label_7[472] = 10'b0000000001;
assign label_7[473] = 10'b0001000000;
assign label_7[474] = 10'b0000000001;
assign label_7[475] = 10'b0000000001;
assign label_7[476] = 10'b0000001000;
assign label_7[477] = 10'b0000100000;
assign label_7[478] = 10'b0000100000;
assign label_7[479] = 10'b0000000001;
assign label_7[480] = 10'b0100000000;
assign label_7[481] = 10'b0100000000;
assign label_7[482] = 10'b0000010000;
assign label_7[483] = 10'b0000010000;
assign label_7[484] = 10'b0001000000;
assign label_7[485] = 10'b0001000000;
assign label_7[486] = 10'b0000010000;
assign label_7[487] = 10'b0000010000;
assign label_7[488] = 10'b0000100000;
assign label_7[489] = 10'b0000100000;
assign label_7[490] = 10'b0001000000;
assign label_7[491] = 10'b0001000000;
assign label_7[492] = 10'b0100000000;
assign label_7[493] = 10'b1000000000;
assign label_7[494] = 10'b0000100000;
assign label_7[495] = 10'b0000000001;
assign label_7[496] = 10'b0000100000;
assign label_7[497] = 10'b0000001000;
assign label_7[498] = 10'b0001000000;
assign label_7[499] = 10'b0000000001;
assign label_7[500] = 10'b0000100000;
assign label_7[501] = 10'b0000100000;
assign label_7[502] = 10'b1000000000;
assign label_7[503] = 10'b0000100000;
assign label_7[504] = 10'b0000000001;
assign label_7[505] = 10'b0001000000;
assign label_7[506] = 10'b0001000000;
assign label_7[507] = 10'b0000000001;
assign label_7[508] = 10'b0000000001;
assign label_7[509] = 10'b0000000001;
assign label_7[510] = 10'b0000000001;
assign label_7[511] = 10'b0000001000;
assign label_7[512] = 10'b0000000010;
assign label_7[513] = 10'b0010000000;
assign label_7[514] = 10'b0000000010;
assign label_7[515] = 10'b0100000000;
assign label_7[516] = 10'b0000000010;
assign label_7[517] = 10'b0001000000;
assign label_7[518] = 10'b0000000100;
assign label_7[519] = 10'b0000000010;
assign label_7[520] = 10'b0000000100;
assign label_7[521] = 10'b0000000010;
assign label_7[522] = 10'b0000001000;
assign label_7[523] = 10'b0000001000;
assign label_7[524] = 10'b0000001000;
assign label_7[525] = 10'b0000001000;
assign label_7[526] = 10'b0000010000;
assign label_7[527] = 10'b0000010000;
assign label_7[528] = 10'b0000100000;
assign label_7[529] = 10'b0000010000;
assign label_7[530] = 10'b0000000100;
assign label_7[531] = 10'b0000000100;
assign label_7[532] = 10'b1000000000;
assign label_7[533] = 10'b0001000000;
assign label_7[534] = 10'b1000000000;
assign label_7[535] = 10'b0000010000;
assign label_7[536] = 10'b0010000000;
assign label_7[537] = 10'b0000000100;
assign label_7[538] = 10'b0000000100;
assign label_7[539] = 10'b0100000000;
assign label_7[540] = 10'b0000000100;
assign label_7[541] = 10'b0000000100;
assign label_7[542] = 10'b0001000000;
assign label_7[543] = 10'b0001000000;
assign label_7[544] = 10'b0000001000;
assign label_7[545] = 10'b0000000010;
assign label_7[546] = 10'b0010000000;
assign label_7[547] = 10'b0001000000;
assign label_7[548] = 10'b0000001000;
assign label_7[549] = 10'b0001000000;
assign label_7[550] = 10'b0000001000;
assign label_7[551] = 10'b0000001000;
assign label_7[552] = 10'b0001000000;
assign label_7[553] = 10'b0100000000;
assign label_7[554] = 10'b0000000100;
assign label_7[555] = 10'b0001000000;
assign label_7[556] = 10'b0001000000;
assign label_7[557] = 10'b0000000100;
assign label_7[558] = 10'b0000000100;
assign label_7[559] = 10'b0000000100;
assign label_7[560] = 10'b0000100000;
assign label_7[561] = 10'b0001000000;
assign label_7[562] = 10'b0000000100;
assign label_7[563] = 10'b0001000000;
assign label_7[564] = 10'b0001000000;
assign label_7[565] = 10'b0100000000;
assign label_7[566] = 10'b0000000100;
assign label_7[567] = 10'b0000000100;
assign label_7[568] = 10'b0000100000;
assign label_7[569] = 10'b0000100000;
assign label_7[570] = 10'b0100000000;
assign label_7[571] = 10'b0000100000;
assign label_7[572] = 10'b0000001000;
assign label_7[573] = 10'b0100000000;
assign label_7[574] = 10'b0000000001;
assign label_7[575] = 10'b0010000000;
assign label_7[576] = 10'b0000000010;
assign label_7[577] = 10'b0000010000;
assign label_7[578] = 10'b0010000000;
assign label_7[579] = 10'b1000000000;
assign label_7[580] = 10'b0000001000;
assign label_7[581] = 10'b0000001000;
assign label_7[582] = 10'b0000000100;
assign label_7[583] = 10'b0001000000;
assign label_7[584] = 10'b0100000000;
assign label_7[585] = 10'b0100000000;
assign label_7[586] = 10'b0000000100;
assign label_7[587] = 10'b0010000000;
assign label_7[588] = 10'b0000000010;
assign label_7[589] = 10'b0100000000;
assign label_7[590] = 10'b0000000100;
assign label_7[591] = 10'b0010000000;
assign label_7[592] = 10'b0000000100;
assign label_7[593] = 10'b0000001000;
assign label_7[594] = 10'b0001000000;
assign label_7[595] = 10'b0000001000;
assign label_7[596] = 10'b0000000100;
assign label_7[597] = 10'b0001000000;
assign label_7[598] = 10'b0000000100;
assign label_7[599] = 10'b0100000000;
assign label_7[600] = 10'b1000000000;
assign label_7[601] = 10'b0100000000;
assign label_7[602] = 10'b0100000000;
assign label_7[603] = 10'b0001000000;
assign label_7[604] = 10'b0001000000;
assign label_7[605] = 10'b0100000000;
assign label_7[606] = 10'b0001000000;
assign label_7[607] = 10'b0000000100;
assign label_7[608] = 10'b0010000000;
assign label_7[609] = 10'b0000001000;
assign label_7[610] = 10'b0000001000;
assign label_7[611] = 10'b0010000000;
assign label_7[612] = 10'b0010000000;
assign label_7[613] = 10'b0010000000;
assign label_7[614] = 10'b0000000100;
assign label_7[615] = 10'b0000001000;
assign label_7[616] = 10'b0000001000;
assign label_7[617] = 10'b0000001000;
assign label_7[618] = 10'b0000001000;
assign label_7[619] = 10'b0000001000;
assign label_7[620] = 10'b0010000000;
assign label_7[621] = 10'b0010000000;
assign label_7[622] = 10'b0010000000;
assign label_7[623] = 10'b0010000000;
assign label_7[624] = 10'b1000000000;
assign label_7[625] = 10'b1000000000;
assign label_7[626] = 10'b1000000000;
assign label_7[627] = 10'b1000000000;
assign label_7[628] = 10'b0010000000;
assign label_7[629] = 10'b0010000000;
assign label_7[630] = 10'b0000001000;
assign label_7[631] = 10'b0000001000;
assign label_7[632] = 10'b0010000000;
assign label_7[633] = 10'b0010000000;
assign label_7[634] = 10'b0100000000;
assign label_7[635] = 10'b0010000000;
assign label_7[636] = 10'b0100000000;
assign label_7[637] = 10'b1000000000;
assign label_7[638] = 10'b0000100000;
assign label_7[639] = 10'b0000001000;
assign label_7[640] = 10'b0000000010;
assign label_7[641] = 10'b0000000010;
assign label_7[642] = 10'b0000100000;
assign label_7[643] = 10'b0000010000;
assign label_7[644] = 10'b0000100000;
assign label_7[645] = 10'b0000010000;
assign label_7[646] = 10'b0001000000;
assign label_7[647] = 10'b0000000100;
assign label_7[648] = 10'b0000010000;
assign label_7[649] = 10'b0001000000;
assign label_7[650] = 10'b0001000000;
assign label_7[651] = 10'b0001000000;
assign label_7[652] = 10'b0000000100;
assign label_7[653] = 10'b0010000000;
assign label_7[654] = 10'b0000010000;
assign label_7[655] = 10'b1000000000;
assign label_7[656] = 10'b0000010000;
assign label_7[657] = 10'b0000010000;
assign label_7[658] = 10'b0001000000;
assign label_7[659] = 10'b0100000000;
assign label_7[660] = 10'b0000000100;
assign label_7[661] = 10'b0001000000;
assign label_7[662] = 10'b0001000000;
assign label_7[663] = 10'b0001000000;
assign label_7[664] = 10'b0000000100;
assign label_7[665] = 10'b1000000000;
assign label_7[666] = 10'b0000000100;
assign label_7[667] = 10'b0000001000;
assign label_7[668] = 10'b0000000100;
assign label_7[669] = 10'b0000000100;
assign label_7[670] = 10'b0000000100;
assign label_7[671] = 10'b0000000100;
assign label_7[672] = 10'b1000000000;
assign label_7[673] = 10'b0001000000;
assign label_7[674] = 10'b0010000000;
assign label_7[675] = 10'b0000001000;
assign label_7[676] = 10'b0010000000;
assign label_7[677] = 10'b0000000100;
assign label_7[678] = 10'b0000001000;
assign label_7[679] = 10'b0000000010;
assign label_7[680] = 10'b0000000100;
assign label_7[681] = 10'b1000000000;
assign label_7[682] = 10'b1000000000;
assign label_7[683] = 10'b0000001000;
assign label_7[684] = 10'b0000100000;
assign label_7[685] = 10'b0100000000;
assign label_7[686] = 10'b0000001000;
assign label_7[687] = 10'b0000001000;
assign label_7[688] = 10'b0010000000;
assign label_7[689] = 10'b1000000000;
assign label_7[690] = 10'b0010000000;
assign label_7[691] = 10'b0000000100;
assign label_7[692] = 10'b0000001000;
assign label_7[693] = 10'b1000000000;
assign label_7[694] = 10'b0000000100;
assign label_7[695] = 10'b0000000100;
assign label_7[696] = 10'b1000000000;
assign label_7[697] = 10'b1000000000;
assign label_7[698] = 10'b0000100000;
assign label_7[699] = 10'b1000000000;
assign label_7[700] = 10'b0100000000;
assign label_7[701] = 10'b1000000000;
assign label_7[702] = 10'b0001000000;
assign label_7[703] = 10'b0000000100;
assign label_7[704] = 10'b0000000100;
assign label_7[705] = 10'b0000100000;
assign label_7[706] = 10'b0000000100;
assign label_7[707] = 10'b0000010000;
assign label_7[708] = 10'b0000000010;
assign label_7[709] = 10'b0001000000;
assign label_7[710] = 10'b0000000010;
assign label_7[711] = 10'b0001000000;
assign label_7[712] = 10'b0000000100;
assign label_7[713] = 10'b0000000100;
assign label_7[714] = 10'b0000000100;
assign label_7[715] = 10'b0000000100;
assign label_7[716] = 10'b0000000001;
assign label_7[717] = 10'b0000000100;
assign label_7[718] = 10'b1000000000;
assign label_7[719] = 10'b1000000000;
assign label_7[720] = 10'b0000000100;
assign label_7[721] = 10'b0100000000;
assign label_7[722] = 10'b0000000100;
assign label_7[723] = 10'b0001000000;
assign label_7[724] = 10'b0000000100;
assign label_7[725] = 10'b0000000100;
assign label_7[726] = 10'b0000000100;
assign label_7[727] = 10'b0001000000;
assign label_7[728] = 10'b0000000100;
assign label_7[729] = 10'b0001000000;
assign label_7[730] = 10'b0001000000;
assign label_7[731] = 10'b0001000000;
assign label_7[732] = 10'b0000000100;
assign label_7[733] = 10'b0000000100;
assign label_7[734] = 10'b1000000000;
assign label_7[735] = 10'b0000010000;
assign label_7[736] = 10'b0100000000;
assign label_7[737] = 10'b0000010000;
assign label_7[738] = 10'b0000010000;
assign label_7[739] = 10'b0000100000;
assign label_7[740] = 10'b0000000010;
assign label_7[741] = 10'b0100000000;
assign label_7[742] = 10'b0000100000;
assign label_7[743] = 10'b0010000000;
assign label_7[744] = 10'b0000001000;
assign label_7[745] = 10'b0100000000;
assign label_7[746] = 10'b0100000000;
assign label_7[747] = 10'b0000000001;
assign label_7[748] = 10'b0010000000;
assign label_7[749] = 10'b0000001000;
assign label_7[750] = 10'b0100000000;
assign label_7[751] = 10'b0000100000;
assign label_7[752] = 10'b0000000100;
assign label_7[753] = 10'b0100000000;
assign label_7[754] = 10'b0000001000;
assign label_7[755] = 10'b0000001000;
assign label_7[756] = 10'b0000000100;
assign label_7[757] = 10'b0100000000;
assign label_7[758] = 10'b0000000100;
assign label_7[759] = 10'b0100000000;
assign label_7[760] = 10'b0100000000;
assign label_7[761] = 10'b0000001000;
assign label_7[762] = 10'b0100000000;
assign label_7[763] = 10'b0000000100;
assign label_7[764] = 10'b0000000100;
assign label_7[765] = 10'b0000000100;
assign label_7[766] = 10'b0000001000;
assign label_7[767] = 10'b1000000000;
assign label_7[768] = 10'b0000100000;
assign label_7[769] = 10'b0000010000;
assign label_7[770] = 10'b0000010000;
assign label_7[771] = 10'b0100000000;
assign label_7[772] = 10'b0100000000;
assign label_7[773] = 10'b0001000000;
assign label_7[774] = 10'b0000100000;
assign label_7[775] = 10'b0000010000;
assign label_7[776] = 10'b0000100000;
assign label_7[777] = 10'b0000001000;
assign label_7[778] = 10'b0001000000;
assign label_7[779] = 10'b0001000000;
assign label_7[780] = 10'b0100000000;
assign label_7[781] = 10'b0100000000;
assign label_7[782] = 10'b0001000000;
assign label_7[783] = 10'b0001000000;
assign label_7[784] = 10'b0000001000;
assign label_7[785] = 10'b0100000000;
assign label_7[786] = 10'b0000100000;
assign label_7[787] = 10'b0000000100;
assign label_7[788] = 10'b0001000000;
assign label_7[789] = 10'b0000000001;
assign label_7[790] = 10'b0001000000;
assign label_7[791] = 10'b0001000000;
assign label_7[792] = 10'b0001000000;
assign label_7[793] = 10'b0100000000;
assign label_7[794] = 10'b0000000100;
assign label_7[795] = 10'b0000000100;
assign label_7[796] = 10'b0001000000;
assign label_7[797] = 10'b0000000001;
assign label_7[798] = 10'b0000000100;
assign label_7[799] = 10'b0100000000;
assign label_7[800] = 10'b0000010000;
assign label_7[801] = 10'b1000000000;
assign label_7[802] = 10'b0000010000;
assign label_7[803] = 10'b0010000000;
assign label_7[804] = 10'b0000010000;
assign label_7[805] = 10'b0000010000;
assign label_7[806] = 10'b0000010000;
assign label_7[807] = 10'b1000000000;
assign label_7[808] = 10'b0000010000;
assign label_7[809] = 10'b0001000000;
assign label_7[810] = 10'b0000010000;
assign label_7[811] = 10'b0100000000;
assign label_7[812] = 10'b0001000000;
assign label_7[813] = 10'b0100000000;
assign label_7[814] = 10'b0000000100;
assign label_7[815] = 10'b0000010000;
assign label_7[816] = 10'b0000010000;
assign label_7[817] = 10'b0001000000;
assign label_7[818] = 10'b0001000000;
assign label_7[819] = 10'b0001000000;
assign label_7[820] = 10'b0000010000;
assign label_7[821] = 10'b0000010000;
assign label_7[822] = 10'b0000001000;
assign label_7[823] = 10'b0000001000;
assign label_7[824] = 10'b0100000000;
assign label_7[825] = 10'b0100000000;
assign label_7[826] = 10'b0100000000;
assign label_7[827] = 10'b0100000000;
assign label_7[828] = 10'b0001000000;
assign label_7[829] = 10'b0001000000;
assign label_7[830] = 10'b0000000100;
assign label_7[831] = 10'b0000000100;
assign label_7[832] = 10'b0000000010;
assign label_7[833] = 10'b0000100000;
assign label_7[834] = 10'b0000010000;
assign label_7[835] = 10'b0100000000;
assign label_7[836] = 10'b0000100000;
assign label_7[837] = 10'b0000001000;
assign label_7[838] = 10'b0100000000;
assign label_7[839] = 10'b0100000000;
assign label_7[840] = 10'b0100000000;
assign label_7[841] = 10'b0100000000;
assign label_7[842] = 10'b0000100000;
assign label_7[843] = 10'b0100000000;
assign label_7[844] = 10'b0000010000;
assign label_7[845] = 10'b0001000000;
assign label_7[846] = 10'b0100000000;
assign label_7[847] = 10'b0100000000;
assign label_7[848] = 10'b0001000000;
assign label_7[849] = 10'b0001000000;
assign label_7[850] = 10'b0000000100;
assign label_7[851] = 10'b0000000100;
assign label_7[852] = 10'b0000000100;
assign label_7[853] = 10'b0000000100;
assign label_7[854] = 10'b0100000000;
assign label_7[855] = 10'b0100000000;
assign label_7[856] = 10'b0001000000;
assign label_7[857] = 10'b0100000000;
assign label_7[858] = 10'b0000000100;
assign label_7[859] = 10'b0001000000;
assign label_7[860] = 10'b0000000100;
assign label_7[861] = 10'b0000000100;
assign label_7[862] = 10'b0000001000;
assign label_7[863] = 10'b0000000100;
assign label_7[864] = 10'b0100000000;
assign label_7[865] = 10'b0000000100;
assign label_7[866] = 10'b0000000010;
assign label_7[867] = 10'b0000100000;
assign label_7[868] = 10'b0001000000;
assign label_7[869] = 10'b0001000000;
assign label_7[870] = 10'b0100000000;
assign label_7[871] = 10'b0000100000;
assign label_7[872] = 10'b0001000000;
assign label_7[873] = 10'b0000000100;
assign label_7[874] = 10'b0000000100;
assign label_7[875] = 10'b0000000100;
assign label_7[876] = 10'b0000000010;
assign label_7[877] = 10'b0000000010;
assign label_7[878] = 10'b0000000010;
assign label_7[879] = 10'b0000000010;
assign label_7[880] = 10'b0000001000;
assign label_7[881] = 10'b0000001000;
assign label_7[882] = 10'b0100000000;
assign label_7[883] = 10'b0001000000;
assign label_7[884] = 10'b0000000100;
assign label_7[885] = 10'b0000000100;
assign label_7[886] = 10'b0000000100;
assign label_7[887] = 10'b0000000100;
assign label_7[888] = 10'b0001000000;
assign label_7[889] = 10'b0001000000;
assign label_7[890] = 10'b0000001000;
assign label_7[891] = 10'b0000001000;
assign label_7[892] = 10'b0001000000;
assign label_7[893] = 10'b0001000000;
assign label_7[894] = 10'b0000000100;
assign label_7[895] = 10'b0000000100;
assign label_7[896] = 10'b0000100000;
assign label_7[897] = 10'b0000100000;
assign label_7[898] = 10'b0000100000;
assign label_7[899] = 10'b0000100000;
assign label_7[900] = 10'b0100000000;
assign label_7[901] = 10'b0100000000;
assign label_7[902] = 10'b0100000000;
assign label_7[903] = 10'b0100000000;
assign label_7[904] = 10'b0001000000;
assign label_7[905] = 10'b0001000000;
assign label_7[906] = 10'b0001000000;
assign label_7[907] = 10'b0001000000;
assign label_7[908] = 10'b0001000000;
assign label_7[909] = 10'b0001000000;
assign label_7[910] = 10'b0001000000;
assign label_7[911] = 10'b0001000000;
assign label_7[912] = 10'b0100000000;
assign label_7[913] = 10'b0100000000;
assign label_7[914] = 10'b0100000000;
assign label_7[915] = 10'b0100000000;
assign label_7[916] = 10'b0000010000;
assign label_7[917] = 10'b0000010000;
assign label_7[918] = 10'b0000010000;
assign label_7[919] = 10'b0000010000;
assign label_7[920] = 10'b0100000000;
assign label_7[921] = 10'b0100000000;
assign label_7[922] = 10'b0100000000;
assign label_7[923] = 10'b0100000000;
assign label_7[924] = 10'b0001000000;
assign label_7[925] = 10'b0001000000;
assign label_7[926] = 10'b0001000000;
assign label_7[927] = 10'b0001000000;
assign label_7[928] = 10'b0001000000;
assign label_7[929] = 10'b0001000000;
assign label_7[930] = 10'b0001000000;
assign label_7[931] = 10'b0001000000;
assign label_7[932] = 10'b0001000000;
assign label_7[933] = 10'b0001000000;
assign label_7[934] = 10'b0001000000;
assign label_7[935] = 10'b0001000000;
assign label_7[936] = 10'b0000000100;
assign label_7[937] = 10'b0000000100;
assign label_7[938] = 10'b0000000100;
assign label_7[939] = 10'b0000000100;
assign label_7[940] = 10'b0001000000;
assign label_7[941] = 10'b0001000000;
assign label_7[942] = 10'b0001000000;
assign label_7[943] = 10'b0001000000;
assign label_7[944] = 10'b0000000100;
assign label_7[945] = 10'b0000000100;
assign label_7[946] = 10'b0000000100;
assign label_7[947] = 10'b0000000100;
assign label_7[948] = 10'b0000000100;
assign label_7[949] = 10'b0000000100;
assign label_7[950] = 10'b0000000100;
assign label_7[951] = 10'b0000000100;
assign label_7[952] = 10'b0000000100;
assign label_7[953] = 10'b0000000100;
assign label_7[954] = 10'b0000000100;
assign label_7[955] = 10'b0000000100;
assign label_7[956] = 10'b0000000100;
assign label_7[957] = 10'b0000000100;
assign label_7[958] = 10'b0000000100;
assign label_7[959] = 10'b0000000100;
assign label_7[960] = 10'b0001000000;
assign label_7[961] = 10'b0001000000;
assign label_7[962] = 10'b0001000000;
assign label_7[963] = 10'b0001000000;
assign label_7[964] = 10'b0000100000;
assign label_7[965] = 10'b0000100000;
assign label_7[966] = 10'b0000100000;
assign label_7[967] = 10'b0000100000;
assign label_7[968] = 10'b0001000000;
assign label_7[969] = 10'b0001000000;
assign label_7[970] = 10'b0001000000;
assign label_7[971] = 10'b0001000000;
assign label_7[972] = 10'b0001000000;
assign label_7[973] = 10'b0001000000;
assign label_7[974] = 10'b0001000000;
assign label_7[975] = 10'b0001000000;
assign label_7[976] = 10'b0000000100;
assign label_7[977] = 10'b0000000100;
assign label_7[978] = 10'b0000000100;
assign label_7[979] = 10'b0000000100;
assign label_7[980] = 10'b0001000000;
assign label_7[981] = 10'b0001000000;
assign label_7[982] = 10'b0001000000;
assign label_7[983] = 10'b0001000000;
assign label_7[984] = 10'b0000000100;
assign label_7[985] = 10'b0000000100;
assign label_7[986] = 10'b0000000100;
assign label_7[987] = 10'b0000000100;
assign label_7[988] = 10'b0000000100;
assign label_7[989] = 10'b0000000100;
assign label_7[990] = 10'b0000000100;
assign label_7[991] = 10'b0000000100;
assign label_7[992] = 10'b0000000010;
assign label_7[993] = 10'b0000000010;
assign label_7[994] = 10'b0000000100;
assign label_7[995] = 10'b0001000000;
assign label_7[996] = 10'b0001000000;
assign label_7[997] = 10'b0001000000;
assign label_7[998] = 10'b0001000000;
assign label_7[999] = 10'b0001000000;
assign label_7[1000] = 10'b0001000000;
assign label_7[1001] = 10'b0000000100;
assign label_7[1002] = 10'b0001000000;
assign label_7[1003] = 10'b0001000000;
assign label_7[1004] = 10'b0001000000;
assign label_7[1005] = 10'b0001000000;
assign label_7[1006] = 10'b0001000000;
assign label_7[1007] = 10'b0001000000;
assign label_7[1008] = 10'b0000000100;
assign label_7[1009] = 10'b0000000100;
assign label_7[1010] = 10'b0000000100;
assign label_7[1011] = 10'b0000000100;
assign label_7[1012] = 10'b0000000100;
assign label_7[1013] = 10'b0000000100;
assign label_7[1014] = 10'b0000000100;
assign label_7[1015] = 10'b0000000100;
assign label_7[1016] = 10'b0000100000;
assign label_7[1017] = 10'b0000100000;
assign label_7[1018] = 10'b0000100000;
assign label_7[1019] = 10'b0000100000;
assign label_7[1020] = 10'b0001000000;
assign label_7[1021] = 10'b0001000000;
assign label_7[1022] = 10'b0000001000;
assign label_7[1023] = 10'b0000001000;
assign label_8[0] = 10'b0010000000;
assign label_8[1] = 10'b0001000000;
assign label_8[2] = 10'b0000010000;
assign label_8[3] = 10'b1000000000;
assign label_8[4] = 10'b0010000000;
assign label_8[5] = 10'b0000100000;
assign label_8[6] = 10'b0010000000;
assign label_8[7] = 10'b1000000000;
assign label_8[8] = 10'b0001000000;
assign label_8[9] = 10'b0000000001;
assign label_8[10] = 10'b0000100000;
assign label_8[11] = 10'b0000010000;
assign label_8[12] = 10'b0001000000;
assign label_8[13] = 10'b0000000001;
assign label_8[14] = 10'b0000000100;
assign label_8[15] = 10'b0000100000;
assign label_8[16] = 10'b0000000010;
assign label_8[17] = 10'b0000001000;
assign label_8[18] = 10'b0000000100;
assign label_8[19] = 10'b0000001000;
assign label_8[20] = 10'b0000000100;
assign label_8[21] = 10'b0100000000;
assign label_8[22] = 10'b0000000100;
assign label_8[23] = 10'b0000001000;
assign label_8[24] = 10'b0000000001;
assign label_8[25] = 10'b0000000001;
assign label_8[26] = 10'b0000000100;
assign label_8[27] = 10'b0000010000;
assign label_8[28] = 10'b0000000100;
assign label_8[29] = 10'b0000000100;
assign label_8[30] = 10'b0000010000;
assign label_8[31] = 10'b0001000000;
assign label_8[32] = 10'b0000000010;
assign label_8[33] = 10'b0000000010;
assign label_8[34] = 10'b0000000100;
assign label_8[35] = 10'b0100000000;
assign label_8[36] = 10'b0010000000;
assign label_8[37] = 10'b0000000100;
assign label_8[38] = 10'b0000000100;
assign label_8[39] = 10'b0000001000;
assign label_8[40] = 10'b0000001000;
assign label_8[41] = 10'b0000100000;
assign label_8[42] = 10'b0000001000;
assign label_8[43] = 10'b0010000000;
assign label_8[44] = 10'b0010000000;
assign label_8[45] = 10'b0000000100;
assign label_8[46] = 10'b0001000000;
assign label_8[47] = 10'b0000000010;
assign label_8[48] = 10'b0000010000;
assign label_8[49] = 10'b0000100000;
assign label_8[50] = 10'b0000001000;
assign label_8[51] = 10'b0000001000;
assign label_8[52] = 10'b0000010000;
assign label_8[53] = 10'b1000000000;
assign label_8[54] = 10'b1000000000;
assign label_8[55] = 10'b0000100000;
assign label_8[56] = 10'b0000000010;
assign label_8[57] = 10'b0000100000;
assign label_8[58] = 10'b0001000000;
assign label_8[59] = 10'b0001000000;
assign label_8[60] = 10'b0000000100;
assign label_8[61] = 10'b0100000000;
assign label_8[62] = 10'b0000001000;
assign label_8[63] = 10'b0100000000;
assign label_8[64] = 10'b0010000000;
assign label_8[65] = 10'b0000000001;
assign label_8[66] = 10'b0010000000;
assign label_8[67] = 10'b0010000000;
assign label_8[68] = 10'b0000100000;
assign label_8[69] = 10'b0100000000;
assign label_8[70] = 10'b1000000000;
assign label_8[71] = 10'b0010000000;
assign label_8[72] = 10'b0000000010;
assign label_8[73] = 10'b0000000100;
assign label_8[74] = 10'b0000100000;
assign label_8[75] = 10'b0100000000;
assign label_8[76] = 10'b0000100000;
assign label_8[77] = 10'b0000100000;
assign label_8[78] = 10'b0010000000;
assign label_8[79] = 10'b0000000001;
assign label_8[80] = 10'b0010000000;
assign label_8[81] = 10'b0000000100;
assign label_8[82] = 10'b0010000000;
assign label_8[83] = 10'b1000000000;
assign label_8[84] = 10'b0000100000;
assign label_8[85] = 10'b0100000000;
assign label_8[86] = 10'b0000000100;
assign label_8[87] = 10'b0000000100;
assign label_8[88] = 10'b1000000000;
assign label_8[89] = 10'b0010000000;
assign label_8[90] = 10'b1000000000;
assign label_8[91] = 10'b0100000000;
assign label_8[92] = 10'b0000100000;
assign label_8[93] = 10'b0000001000;
assign label_8[94] = 10'b0100000000;
assign label_8[95] = 10'b0100000000;
assign label_8[96] = 10'b0000000010;
assign label_8[97] = 10'b0001000000;
assign label_8[98] = 10'b1000000000;
assign label_8[99] = 10'b0001000000;
assign label_8[100] = 10'b0010000000;
assign label_8[101] = 10'b0100000000;
assign label_8[102] = 10'b0000000010;
assign label_8[103] = 10'b1000000000;
assign label_8[104] = 10'b0010000000;
assign label_8[105] = 10'b0010000000;
assign label_8[106] = 10'b0000000001;
assign label_8[107] = 10'b0000000001;
assign label_8[108] = 10'b1000000000;
assign label_8[109] = 10'b0100000000;
assign label_8[110] = 10'b0100000000;
assign label_8[111] = 10'b0100000000;
assign label_8[112] = 10'b0010000000;
assign label_8[113] = 10'b0010000000;
assign label_8[114] = 10'b0100000000;
assign label_8[115] = 10'b0000001000;
assign label_8[116] = 10'b0000000001;
assign label_8[117] = 10'b0000000001;
assign label_8[118] = 10'b0100000000;
assign label_8[119] = 10'b0100000000;
assign label_8[120] = 10'b0100000000;
assign label_8[121] = 10'b0000000100;
assign label_8[122] = 10'b0000000001;
assign label_8[123] = 10'b0001000000;
assign label_8[124] = 10'b0100000000;
assign label_8[125] = 10'b0100000000;
assign label_8[126] = 10'b0000001000;
assign label_8[127] = 10'b0100000000;
assign label_8[128] = 10'b0010000000;
assign label_8[129] = 10'b0001000000;
assign label_8[130] = 10'b0000001000;
assign label_8[131] = 10'b0000000100;
assign label_8[132] = 10'b0000001000;
assign label_8[133] = 10'b0100000000;
assign label_8[134] = 10'b0000000100;
assign label_8[135] = 10'b0000001000;
assign label_8[136] = 10'b0010000000;
assign label_8[137] = 10'b0000001000;
assign label_8[138] = 10'b0000001000;
assign label_8[139] = 10'b0000100000;
assign label_8[140] = 10'b0010000000;
assign label_8[141] = 10'b0000000010;
assign label_8[142] = 10'b0000001000;
assign label_8[143] = 10'b0000000001;
assign label_8[144] = 10'b0010000000;
assign label_8[145] = 10'b0000000100;
assign label_8[146] = 10'b0000000100;
assign label_8[147] = 10'b0000000001;
assign label_8[148] = 10'b0000001000;
assign label_8[149] = 10'b0000100000;
assign label_8[150] = 10'b0000001000;
assign label_8[151] = 10'b0000001000;
assign label_8[152] = 10'b0000001000;
assign label_8[153] = 10'b0010000000;
assign label_8[154] = 10'b0000100000;
assign label_8[155] = 10'b0000001000;
assign label_8[156] = 10'b0001000000;
assign label_8[157] = 10'b0000001000;
assign label_8[158] = 10'b0100000000;
assign label_8[159] = 10'b0000000100;
assign label_8[160] = 10'b0010000000;
assign label_8[161] = 10'b1000000000;
assign label_8[162] = 10'b0010000000;
assign label_8[163] = 10'b1000000000;
assign label_8[164] = 10'b0000000001;
assign label_8[165] = 10'b0010000000;
assign label_8[166] = 10'b0000000001;
assign label_8[167] = 10'b0000000100;
assign label_8[168] = 10'b0000010000;
assign label_8[169] = 10'b1000000000;
assign label_8[170] = 10'b1000000000;
assign label_8[171] = 10'b0000100000;
assign label_8[172] = 10'b0000100000;
assign label_8[173] = 10'b0000001000;
assign label_8[174] = 10'b0000010000;
assign label_8[175] = 10'b1000000000;
assign label_8[176] = 10'b0010000000;
assign label_8[177] = 10'b0010000000;
assign label_8[178] = 10'b0001000000;
assign label_8[179] = 10'b0001000000;
assign label_8[180] = 10'b1000000000;
assign label_8[181] = 10'b0000000001;
assign label_8[182] = 10'b1000000000;
assign label_8[183] = 10'b1000000000;
assign label_8[184] = 10'b0000000001;
assign label_8[185] = 10'b0001000000;
assign label_8[186] = 10'b0001000000;
assign label_8[187] = 10'b0001000000;
assign label_8[188] = 10'b0000000001;
assign label_8[189] = 10'b0000000001;
assign label_8[190] = 10'b0000000001;
assign label_8[191] = 10'b0001000000;
assign label_8[192] = 10'b0000001000;
assign label_8[193] = 10'b0000000010;
assign label_8[194] = 10'b0000001000;
assign label_8[195] = 10'b0000001000;
assign label_8[196] = 10'b0000010000;
assign label_8[197] = 10'b0000001000;
assign label_8[198] = 10'b0000010000;
assign label_8[199] = 10'b1000000000;
assign label_8[200] = 10'b0100000000;
assign label_8[201] = 10'b0000000100;
assign label_8[202] = 10'b0000000100;
assign label_8[203] = 10'b0000000100;
assign label_8[204] = 10'b0001000000;
assign label_8[205] = 10'b0100000000;
assign label_8[206] = 10'b0100000000;
assign label_8[207] = 10'b0000000100;
assign label_8[208] = 10'b0000100000;
assign label_8[209] = 10'b0000100000;
assign label_8[210] = 10'b0000100000;
assign label_8[211] = 10'b0000100000;
assign label_8[212] = 10'b0000001000;
assign label_8[213] = 10'b0000001000;
assign label_8[214] = 10'b0100000000;
assign label_8[215] = 10'b0100000000;
assign label_8[216] = 10'b0010000000;
assign label_8[217] = 10'b0000001000;
assign label_8[218] = 10'b0000001000;
assign label_8[219] = 10'b0000001000;
assign label_8[220] = 10'b0000100000;
assign label_8[221] = 10'b0000000100;
assign label_8[222] = 10'b0100000000;
assign label_8[223] = 10'b0000001000;
assign label_8[224] = 10'b0000000100;
assign label_8[225] = 10'b0000000100;
assign label_8[226] = 10'b0001000000;
assign label_8[227] = 10'b0000000100;
assign label_8[228] = 10'b0000000100;
assign label_8[229] = 10'b0000001000;
assign label_8[230] = 10'b0001000000;
assign label_8[231] = 10'b0001000000;
assign label_8[232] = 10'b0000100000;
assign label_8[233] = 10'b0001000000;
assign label_8[234] = 10'b0000000100;
assign label_8[235] = 10'b0000000100;
assign label_8[236] = 10'b0000100000;
assign label_8[237] = 10'b0001000000;
assign label_8[238] = 10'b0000001000;
assign label_8[239] = 10'b0000000100;
assign label_8[240] = 10'b0000001000;
assign label_8[241] = 10'b0000000100;
assign label_8[242] = 10'b0100000000;
assign label_8[243] = 10'b0000001000;
assign label_8[244] = 10'b0000001000;
assign label_8[245] = 10'b0100000000;
assign label_8[246] = 10'b0000001000;
assign label_8[247] = 10'b0000000100;
assign label_8[248] = 10'b0000001000;
assign label_8[249] = 10'b0000100000;
assign label_8[250] = 10'b0100000000;
assign label_8[251] = 10'b0000000100;
assign label_8[252] = 10'b0001000000;
assign label_8[253] = 10'b0000000001;
assign label_8[254] = 10'b0000001000;
assign label_8[255] = 10'b0000001000;
assign label_8[256] = 10'b0000010000;
assign label_8[257] = 10'b0000010000;
assign label_8[258] = 10'b0010000000;
assign label_8[259] = 10'b1000000000;
assign label_8[260] = 10'b0000010000;
assign label_8[261] = 10'b0000010000;
assign label_8[262] = 10'b0010000000;
assign label_8[263] = 10'b1000000000;
assign label_8[264] = 10'b0000100000;
assign label_8[265] = 10'b0000000010;
assign label_8[266] = 10'b0000000010;
assign label_8[267] = 10'b0000001000;
assign label_8[268] = 10'b0010000000;
assign label_8[269] = 10'b0000010000;
assign label_8[270] = 10'b0010000000;
assign label_8[271] = 10'b0010000000;
assign label_8[272] = 10'b0000100000;
assign label_8[273] = 10'b0000001000;
assign label_8[274] = 10'b0000000100;
assign label_8[275] = 10'b0000000001;
assign label_8[276] = 10'b0000001000;
assign label_8[277] = 10'b0000100000;
assign label_8[278] = 10'b0000000001;
assign label_8[279] = 10'b0000000001;
assign label_8[280] = 10'b0000100000;
assign label_8[281] = 10'b0000100000;
assign label_8[282] = 10'b0000001000;
assign label_8[283] = 10'b0100000000;
assign label_8[284] = 10'b0000100000;
assign label_8[285] = 10'b0000100000;
assign label_8[286] = 10'b0000000100;
assign label_8[287] = 10'b0000000001;
assign label_8[288] = 10'b1000000000;
assign label_8[289] = 10'b0000100000;
assign label_8[290] = 10'b1000000000;
assign label_8[291] = 10'b0000100000;
assign label_8[292] = 10'b0010000000;
assign label_8[293] = 10'b1000000000;
assign label_8[294] = 10'b1000000000;
assign label_8[295] = 10'b0100000000;
assign label_8[296] = 10'b0000100000;
assign label_8[297] = 10'b0100000000;
assign label_8[298] = 10'b0100000000;
assign label_8[299] = 10'b0100000000;
assign label_8[300] = 10'b0000001000;
assign label_8[301] = 10'b0000001000;
assign label_8[302] = 10'b0000001000;
assign label_8[303] = 10'b0000000001;
assign label_8[304] = 10'b0000100000;
assign label_8[305] = 10'b0000000001;
assign label_8[306] = 10'b0000100000;
assign label_8[307] = 10'b0100000000;
assign label_8[308] = 10'b0000100000;
assign label_8[309] = 10'b0000000001;
assign label_8[310] = 10'b0000000100;
assign label_8[311] = 10'b0100000000;
assign label_8[312] = 10'b0000001000;
assign label_8[313] = 10'b0000000100;
assign label_8[314] = 10'b0000001000;
assign label_8[315] = 10'b0000001000;
assign label_8[316] = 10'b0000001000;
assign label_8[317] = 10'b0000100000;
assign label_8[318] = 10'b0000100000;
assign label_8[319] = 10'b0000001000;
assign label_8[320] = 10'b0010000000;
assign label_8[321] = 10'b0000000001;
assign label_8[322] = 10'b0000000100;
assign label_8[323] = 10'b0000000001;
assign label_8[324] = 10'b0001000000;
assign label_8[325] = 10'b0000001000;
assign label_8[326] = 10'b0000100000;
assign label_8[327] = 10'b0100000000;
assign label_8[328] = 10'b0000000100;
assign label_8[329] = 10'b0000000001;
assign label_8[330] = 10'b0000000001;
assign label_8[331] = 10'b0000000001;
assign label_8[332] = 10'b0000100000;
assign label_8[333] = 10'b0000000100;
assign label_8[334] = 10'b0000000001;
assign label_8[335] = 10'b0000000100;
assign label_8[336] = 10'b0000100000;
assign label_8[337] = 10'b0000100000;
assign label_8[338] = 10'b0000001000;
assign label_8[339] = 10'b0000001000;
assign label_8[340] = 10'b0000010000;
assign label_8[341] = 10'b0100000000;
assign label_8[342] = 10'b0000100000;
assign label_8[343] = 10'b0000000001;
assign label_8[344] = 10'b0010000000;
assign label_8[345] = 10'b0000001000;
assign label_8[346] = 10'b0010000000;
assign label_8[347] = 10'b0010000000;
assign label_8[348] = 10'b0000001000;
assign label_8[349] = 10'b0000000001;
assign label_8[350] = 10'b0000001000;
assign label_8[351] = 10'b0000000001;
assign label_8[352] = 10'b0000001000;
assign label_8[353] = 10'b0000001000;
assign label_8[354] = 10'b0000001000;
assign label_8[355] = 10'b0000001000;
assign label_8[356] = 10'b0000001000;
assign label_8[357] = 10'b0000001000;
assign label_8[358] = 10'b0100000000;
assign label_8[359] = 10'b0000001000;
assign label_8[360] = 10'b0000000100;
assign label_8[361] = 10'b0000000100;
assign label_8[362] = 10'b0000000100;
assign label_8[363] = 10'b0000000100;
assign label_8[364] = 10'b0000001000;
assign label_8[365] = 10'b0000001000;
assign label_8[366] = 10'b0000100000;
assign label_8[367] = 10'b0000100000;
assign label_8[368] = 10'b0000001000;
assign label_8[369] = 10'b0000100000;
assign label_8[370] = 10'b0000100000;
assign label_8[371] = 10'b0000100000;
assign label_8[372] = 10'b0000100000;
assign label_8[373] = 10'b0000000100;
assign label_8[374] = 10'b0000001000;
assign label_8[375] = 10'b0000001000;
assign label_8[376] = 10'b0000100000;
assign label_8[377] = 10'b0000010000;
assign label_8[378] = 10'b0000100000;
assign label_8[379] = 10'b0000001000;
assign label_8[380] = 10'b0000100000;
assign label_8[381] = 10'b0000100000;
assign label_8[382] = 10'b0000100000;
assign label_8[383] = 10'b0000100000;
assign label_8[384] = 10'b0000010000;
assign label_8[385] = 10'b0001000000;
assign label_8[386] = 10'b1000000000;
assign label_8[387] = 10'b0000100000;
assign label_8[388] = 10'b1000000000;
assign label_8[389] = 10'b0000010000;
assign label_8[390] = 10'b0000010000;
assign label_8[391] = 10'b0000010000;
assign label_8[392] = 10'b0001000000;
assign label_8[393] = 10'b0100000000;
assign label_8[394] = 10'b0000100000;
assign label_8[395] = 10'b0100000000;
assign label_8[396] = 10'b0100000000;
assign label_8[397] = 10'b0000100000;
assign label_8[398] = 10'b0000010000;
assign label_8[399] = 10'b0100000000;
assign label_8[400] = 10'b1000000000;
assign label_8[401] = 10'b0000001000;
assign label_8[402] = 10'b0100000000;
assign label_8[403] = 10'b1000000000;
assign label_8[404] = 10'b0000100000;
assign label_8[405] = 10'b0000001000;
assign label_8[406] = 10'b1000000000;
assign label_8[407] = 10'b0000001000;
assign label_8[408] = 10'b0000010000;
assign label_8[409] = 10'b0100000000;
assign label_8[410] = 10'b0000010000;
assign label_8[411] = 10'b0100000000;
assign label_8[412] = 10'b0001000000;
assign label_8[413] = 10'b0000100000;
assign label_8[414] = 10'b0100000000;
assign label_8[415] = 10'b0000001000;
assign label_8[416] = 10'b0000100000;
assign label_8[417] = 10'b0000000001;
assign label_8[418] = 10'b0000100000;
assign label_8[419] = 10'b0000001000;
assign label_8[420] = 10'b0000100000;
assign label_8[421] = 10'b1000000000;
assign label_8[422] = 10'b0000010000;
assign label_8[423] = 10'b0100000000;
assign label_8[424] = 10'b0000001000;
assign label_8[425] = 10'b0000100000;
assign label_8[426] = 10'b0000100000;
assign label_8[427] = 10'b0000100000;
assign label_8[428] = 10'b0000001000;
assign label_8[429] = 10'b0000001000;
assign label_8[430] = 10'b0000100000;
assign label_8[431] = 10'b0000001000;
assign label_8[432] = 10'b0000100000;
assign label_8[433] = 10'b0000100000;
assign label_8[434] = 10'b0100000000;
assign label_8[435] = 10'b0000100000;
assign label_8[436] = 10'b1000000000;
assign label_8[437] = 10'b0000001000;
assign label_8[438] = 10'b0000100000;
assign label_8[439] = 10'b0000001000;
assign label_8[440] = 10'b1000000000;
assign label_8[441] = 10'b0000010000;
assign label_8[442] = 10'b0000010000;
assign label_8[443] = 10'b0100000000;
assign label_8[444] = 10'b0000001000;
assign label_8[445] = 10'b0100000000;
assign label_8[446] = 10'b1000000000;
assign label_8[447] = 10'b0000001000;
assign label_8[448] = 10'b0100000000;
assign label_8[449] = 10'b0000000100;
assign label_8[450] = 10'b0100000000;
assign label_8[451] = 10'b0100000000;
assign label_8[452] = 10'b0100000000;
assign label_8[453] = 10'b0100000000;
assign label_8[454] = 10'b0010000000;
assign label_8[455] = 10'b0010000000;
assign label_8[456] = 10'b0100000000;
assign label_8[457] = 10'b0100000000;
assign label_8[458] = 10'b0100000000;
assign label_8[459] = 10'b0000000010;
assign label_8[460] = 10'b0100000000;
assign label_8[461] = 10'b0100000000;
assign label_8[462] = 10'b0100000000;
assign label_8[463] = 10'b0100000000;
assign label_8[464] = 10'b0010000000;
assign label_8[465] = 10'b0100000000;
assign label_8[466] = 10'b0100000000;
assign label_8[467] = 10'b0100000000;
assign label_8[468] = 10'b0010000000;
assign label_8[469] = 10'b0100000000;
assign label_8[470] = 10'b0100000000;
assign label_8[471] = 10'b0100000000;
assign label_8[472] = 10'b0000000100;
assign label_8[473] = 10'b0000000100;
assign label_8[474] = 10'b0000000100;
assign label_8[475] = 10'b0000000100;
assign label_8[476] = 10'b0100000000;
assign label_8[477] = 10'b0000001000;
assign label_8[478] = 10'b0000100000;
assign label_8[479] = 10'b0001000000;
assign label_8[480] = 10'b0000010000;
assign label_8[481] = 10'b0001000000;
assign label_8[482] = 10'b0100000000;
assign label_8[483] = 10'b0100000000;
assign label_8[484] = 10'b0001000000;
assign label_8[485] = 10'b0100000000;
assign label_8[486] = 10'b0001000000;
assign label_8[487] = 10'b0100000000;
assign label_8[488] = 10'b0000100000;
assign label_8[489] = 10'b0000100000;
assign label_8[490] = 10'b0001000000;
assign label_8[491] = 10'b0001000000;
assign label_8[492] = 10'b0000000001;
assign label_8[493] = 10'b0001000000;
assign label_8[494] = 10'b0001000000;
assign label_8[495] = 10'b0000000100;
assign label_8[496] = 10'b0001000000;
assign label_8[497] = 10'b0100000000;
assign label_8[498] = 10'b0000100000;
assign label_8[499] = 10'b0000010000;
assign label_8[500] = 10'b0000000001;
assign label_8[501] = 10'b0000000100;
assign label_8[502] = 10'b0001000000;
assign label_8[503] = 10'b0100000000;
assign label_8[504] = 10'b1000000000;
assign label_8[505] = 10'b0000000001;
assign label_8[506] = 10'b0100000000;
assign label_8[507] = 10'b0100000000;
assign label_8[508] = 10'b0000000001;
assign label_8[509] = 10'b0100000000;
assign label_8[510] = 10'b0100000000;
assign label_8[511] = 10'b0100000000;
assign label_8[512] = 10'b0010000000;
assign label_8[513] = 10'b0000010000;
assign label_8[514] = 10'b0000010000;
assign label_8[515] = 10'b0000010000;
assign label_8[516] = 10'b1000000000;
assign label_8[517] = 10'b0000000100;
assign label_8[518] = 10'b0000000100;
assign label_8[519] = 10'b0000001000;
assign label_8[520] = 10'b0010000000;
assign label_8[521] = 10'b0000100000;
assign label_8[522] = 10'b0010000000;
assign label_8[523] = 10'b1000000000;
assign label_8[524] = 10'b0000010000;
assign label_8[525] = 10'b0000010000;
assign label_8[526] = 10'b0000010000;
assign label_8[527] = 10'b1000000000;
assign label_8[528] = 10'b0000010000;
assign label_8[529] = 10'b0001000000;
assign label_8[530] = 10'b0000100000;
assign label_8[531] = 10'b1000000000;
assign label_8[532] = 10'b0000000100;
assign label_8[533] = 10'b1000000000;
assign label_8[534] = 10'b0000000001;
assign label_8[535] = 10'b0000000001;
assign label_8[536] = 10'b0000000100;
assign label_8[537] = 10'b0001000000;
assign label_8[538] = 10'b0000100000;
assign label_8[539] = 10'b0000100000;
assign label_8[540] = 10'b0000000001;
assign label_8[541] = 10'b0100000000;
assign label_8[542] = 10'b0000000100;
assign label_8[543] = 10'b0000000100;
assign label_8[544] = 10'b0000010000;
assign label_8[545] = 10'b0000010000;
assign label_8[546] = 10'b0000001000;
assign label_8[547] = 10'b0000000100;
assign label_8[548] = 10'b0000000100;
assign label_8[549] = 10'b0000000100;
assign label_8[550] = 10'b0000001000;
assign label_8[551] = 10'b0000001000;
assign label_8[552] = 10'b0000000100;
assign label_8[553] = 10'b0000000100;
assign label_8[554] = 10'b0000000100;
assign label_8[555] = 10'b0000000100;
assign label_8[556] = 10'b0000000100;
assign label_8[557] = 10'b0000000100;
assign label_8[558] = 10'b0000000100;
assign label_8[559] = 10'b0000000100;
assign label_8[560] = 10'b0000010000;
assign label_8[561] = 10'b0000010000;
assign label_8[562] = 10'b0000010000;
assign label_8[563] = 10'b0000010000;
assign label_8[564] = 10'b0001000000;
assign label_8[565] = 10'b1000000000;
assign label_8[566] = 10'b0000010000;
assign label_8[567] = 10'b0000010000;
assign label_8[568] = 10'b0001000000;
assign label_8[569] = 10'b0001000000;
assign label_8[570] = 10'b0001000000;
assign label_8[571] = 10'b0001000000;
assign label_8[572] = 10'b0000010000;
assign label_8[573] = 10'b0000010000;
assign label_8[574] = 10'b0001000000;
assign label_8[575] = 10'b0001000000;
assign label_8[576] = 10'b0000000100;
assign label_8[577] = 10'b0010000000;
assign label_8[578] = 10'b0000000100;
assign label_8[579] = 10'b0000000100;
assign label_8[580] = 10'b0010000000;
assign label_8[581] = 10'b1000000000;
assign label_8[582] = 10'b0100000000;
assign label_8[583] = 10'b0000010000;
assign label_8[584] = 10'b0000010000;
assign label_8[585] = 10'b0000000100;
assign label_8[586] = 10'b0000000100;
assign label_8[587] = 10'b0000010000;
assign label_8[588] = 10'b0000001000;
assign label_8[589] = 10'b0000000100;
assign label_8[590] = 10'b0001000000;
assign label_8[591] = 10'b0100000000;
assign label_8[592] = 10'b1000000000;
assign label_8[593] = 10'b0000100000;
assign label_8[594] = 10'b0000100000;
assign label_8[595] = 10'b1000000000;
assign label_8[596] = 10'b1000000000;
assign label_8[597] = 10'b0001000000;
assign label_8[598] = 10'b1000000000;
assign label_8[599] = 10'b0001000000;
assign label_8[600] = 10'b0000000001;
assign label_8[601] = 10'b0000000001;
assign label_8[602] = 10'b0000010000;
assign label_8[603] = 10'b0000100000;
assign label_8[604] = 10'b0000010000;
assign label_8[605] = 10'b0000010000;
assign label_8[606] = 10'b0000010000;
assign label_8[607] = 10'b1000000000;
assign label_8[608] = 10'b0000000001;
assign label_8[609] = 10'b0000000001;
assign label_8[610] = 10'b0000100000;
assign label_8[611] = 10'b0000100000;
assign label_8[612] = 10'b0000100000;
assign label_8[613] = 10'b0000100000;
assign label_8[614] = 10'b1000000000;
assign label_8[615] = 10'b0010000000;
assign label_8[616] = 10'b0000100000;
assign label_8[617] = 10'b0100000000;
assign label_8[618] = 10'b0000100000;
assign label_8[619] = 10'b0100000000;
assign label_8[620] = 10'b0000001000;
assign label_8[621] = 10'b0100000000;
assign label_8[622] = 10'b0000000001;
assign label_8[623] = 10'b0000000001;
assign label_8[624] = 10'b0000001000;
assign label_8[625] = 10'b0000001000;
assign label_8[626] = 10'b0000100000;
assign label_8[627] = 10'b0000100000;
assign label_8[628] = 10'b0000001000;
assign label_8[629] = 10'b0100000000;
assign label_8[630] = 10'b0000001000;
assign label_8[631] = 10'b0100000000;
assign label_8[632] = 10'b0000001000;
assign label_8[633] = 10'b0100000000;
assign label_8[634] = 10'b0000100000;
assign label_8[635] = 10'b0000100000;
assign label_8[636] = 10'b0000100000;
assign label_8[637] = 10'b0100000000;
assign label_8[638] = 10'b0100000000;
assign label_8[639] = 10'b0100000000;
assign label_8[640] = 10'b0000000001;
assign label_8[641] = 10'b0001000000;
assign label_8[642] = 10'b0000000001;
assign label_8[643] = 10'b0000000001;
assign label_8[644] = 10'b0000000001;
assign label_8[645] = 10'b0000000001;
assign label_8[646] = 10'b0000100000;
assign label_8[647] = 10'b0000000001;
assign label_8[648] = 10'b0000100000;
assign label_8[649] = 10'b0000000001;
assign label_8[650] = 10'b0000000001;
assign label_8[651] = 10'b0000000001;
assign label_8[652] = 10'b0000100000;
assign label_8[653] = 10'b0000000001;
assign label_8[654] = 10'b0000001000;
assign label_8[655] = 10'b0000100000;
assign label_8[656] = 10'b0000100000;
assign label_8[657] = 10'b0001000000;
assign label_8[658] = 10'b0000000100;
assign label_8[659] = 10'b0000000100;
assign label_8[660] = 10'b0000000100;
assign label_8[661] = 10'b0000000100;
assign label_8[662] = 10'b0001000000;
assign label_8[663] = 10'b0000100000;
assign label_8[664] = 10'b0000100000;
assign label_8[665] = 10'b1000000000;
assign label_8[666] = 10'b0000100000;
assign label_8[667] = 10'b0000100000;
assign label_8[668] = 10'b0000100000;
assign label_8[669] = 10'b0001000000;
assign label_8[670] = 10'b0100000000;
assign label_8[671] = 10'b0000000001;
assign label_8[672] = 10'b0010000000;
assign label_8[673] = 10'b0000000001;
assign label_8[674] = 10'b0000010000;
assign label_8[675] = 10'b0000100000;
assign label_8[676] = 10'b0001000000;
assign label_8[677] = 10'b0000000001;
assign label_8[678] = 10'b0001000000;
assign label_8[679] = 10'b0000000001;
assign label_8[680] = 10'b1000000000;
assign label_8[681] = 10'b0000010000;
assign label_8[682] = 10'b0000010000;
assign label_8[683] = 10'b1000000000;
assign label_8[684] = 10'b0000000100;
assign label_8[685] = 10'b0000000100;
assign label_8[686] = 10'b0000100000;
assign label_8[687] = 10'b0001000000;
assign label_8[688] = 10'b0000010000;
assign label_8[689] = 10'b1000000000;
assign label_8[690] = 10'b0001000000;
assign label_8[691] = 10'b0000000100;
assign label_8[692] = 10'b0000010000;
assign label_8[693] = 10'b1000000000;
assign label_8[694] = 10'b0000000100;
assign label_8[695] = 10'b0000000001;
assign label_8[696] = 10'b1000000000;
assign label_8[697] = 10'b0000100000;
assign label_8[698] = 10'b0000010000;
assign label_8[699] = 10'b1000000000;
assign label_8[700] = 10'b0000000001;
assign label_8[701] = 10'b0000000001;
assign label_8[702] = 10'b0001000000;
assign label_8[703] = 10'b0000100000;
assign label_8[704] = 10'b0000010000;
assign label_8[705] = 10'b0000100000;
assign label_8[706] = 10'b0000010000;
assign label_8[707] = 10'b0000010000;
assign label_8[708] = 10'b0000100000;
assign label_8[709] = 10'b0001000000;
assign label_8[710] = 10'b0100000000;
assign label_8[711] = 10'b0000000001;
assign label_8[712] = 10'b0000001000;
assign label_8[713] = 10'b0100000000;
assign label_8[714] = 10'b0000100000;
assign label_8[715] = 10'b0100000000;
assign label_8[716] = 10'b0000100000;
assign label_8[717] = 10'b0100000000;
assign label_8[718] = 10'b0000001000;
assign label_8[719] = 10'b0100000000;
assign label_8[720] = 10'b0000001000;
assign label_8[721] = 10'b0000100000;
assign label_8[722] = 10'b0000100000;
assign label_8[723] = 10'b0000100000;
assign label_8[724] = 10'b0100000000;
assign label_8[725] = 10'b0000100000;
assign label_8[726] = 10'b0100000000;
assign label_8[727] = 10'b0000000001;
assign label_8[728] = 10'b0000010000;
assign label_8[729] = 10'b1000000000;
assign label_8[730] = 10'b1000000000;
assign label_8[731] = 10'b0000010000;
assign label_8[732] = 10'b0000010000;
assign label_8[733] = 10'b0100000000;
assign label_8[734] = 10'b0000100000;
assign label_8[735] = 10'b0100000000;
assign label_8[736] = 10'b0100000000;
assign label_8[737] = 10'b0000000100;
assign label_8[738] = 10'b0000000100;
assign label_8[739] = 10'b0000000100;
assign label_8[740] = 10'b0000000100;
assign label_8[741] = 10'b0100000000;
assign label_8[742] = 10'b0100000000;
assign label_8[743] = 10'b0000001000;
assign label_8[744] = 10'b0001000000;
assign label_8[745] = 10'b0100000000;
assign label_8[746] = 10'b0001000000;
assign label_8[747] = 10'b0100000000;
assign label_8[748] = 10'b0000010000;
assign label_8[749] = 10'b0000000100;
assign label_8[750] = 10'b0000000001;
assign label_8[751] = 10'b0100000000;
assign label_8[752] = 10'b0000000100;
assign label_8[753] = 10'b0000000100;
assign label_8[754] = 10'b0000000001;
assign label_8[755] = 10'b0000000100;
assign label_8[756] = 10'b0000000100;
assign label_8[757] = 10'b0100000000;
assign label_8[758] = 10'b0100000000;
assign label_8[759] = 10'b0001000000;
assign label_8[760] = 10'b0000001000;
assign label_8[761] = 10'b0000001000;
assign label_8[762] = 10'b0100000000;
assign label_8[763] = 10'b0000000100;
assign label_8[764] = 10'b0000000001;
assign label_8[765] = 10'b0000000001;
assign label_8[766] = 10'b0100000000;
assign label_8[767] = 10'b0100000000;
assign label_8[768] = 10'b0000000100;
assign label_8[769] = 10'b0001000000;
assign label_8[770] = 10'b0000000100;
assign label_8[771] = 10'b0000000100;
assign label_8[772] = 10'b0000010000;
assign label_8[773] = 10'b1000000000;
assign label_8[774] = 10'b0000100000;
assign label_8[775] = 10'b0000000100;
assign label_8[776] = 10'b0000000010;
assign label_8[777] = 10'b0000000010;
assign label_8[778] = 10'b0000000010;
assign label_8[779] = 10'b0000000010;
assign label_8[780] = 10'b0100000000;
assign label_8[781] = 10'b0100000000;
assign label_8[782] = 10'b0000010000;
assign label_8[783] = 10'b0000010000;
assign label_8[784] = 10'b0001000000;
assign label_8[785] = 10'b0001000000;
assign label_8[786] = 10'b0001000000;
assign label_8[787] = 10'b0000000100;
assign label_8[788] = 10'b0000010000;
assign label_8[789] = 10'b0000010000;
assign label_8[790] = 10'b0000100000;
assign label_8[791] = 10'b0000100000;
assign label_8[792] = 10'b0000000100;
assign label_8[793] = 10'b0001000000;
assign label_8[794] = 10'b0001000000;
assign label_8[795] = 10'b1000000000;
assign label_8[796] = 10'b0000010000;
assign label_8[797] = 10'b0000000100;
assign label_8[798] = 10'b0000000001;
assign label_8[799] = 10'b0000000100;
assign label_8[800] = 10'b0001000000;
assign label_8[801] = 10'b0000000100;
assign label_8[802] = 10'b0000000100;
assign label_8[803] = 10'b0001000000;
assign label_8[804] = 10'b0100000000;
assign label_8[805] = 10'b0000010000;
assign label_8[806] = 10'b0010000000;
assign label_8[807] = 10'b0010000000;
assign label_8[808] = 10'b0000000100;
assign label_8[809] = 10'b0000000100;
assign label_8[810] = 10'b0000000100;
assign label_8[811] = 10'b0000000100;
assign label_8[812] = 10'b0000000100;
assign label_8[813] = 10'b0000000100;
assign label_8[814] = 10'b0000000100;
assign label_8[815] = 10'b0000000100;
assign label_8[816] = 10'b0001000000;
assign label_8[817] = 10'b0001000000;
assign label_8[818] = 10'b0000000001;
assign label_8[819] = 10'b0000000100;
assign label_8[820] = 10'b0000010000;
assign label_8[821] = 10'b0000010000;
assign label_8[822] = 10'b0000000100;
assign label_8[823] = 10'b0000000001;
assign label_8[824] = 10'b0000000001;
assign label_8[825] = 10'b0000000001;
assign label_8[826] = 10'b0001000000;
assign label_8[827] = 10'b0000000001;
assign label_8[828] = 10'b0000010000;
assign label_8[829] = 10'b0000010000;
assign label_8[830] = 10'b0000000100;
assign label_8[831] = 10'b0000000100;
assign label_8[832] = 10'b0000000100;
assign label_8[833] = 10'b0000000100;
assign label_8[834] = 10'b1000000000;
assign label_8[835] = 10'b0000001000;
assign label_8[836] = 10'b0100000000;
assign label_8[837] = 10'b0000000100;
assign label_8[838] = 10'b0000100000;
assign label_8[839] = 10'b0000100000;
assign label_8[840] = 10'b1000000000;
assign label_8[841] = 10'b1000000000;
assign label_8[842] = 10'b0001000000;
assign label_8[843] = 10'b0000000100;
assign label_8[844] = 10'b0001000000;
assign label_8[845] = 10'b0000100000;
assign label_8[846] = 10'b0000000001;
assign label_8[847] = 10'b0000000001;
assign label_8[848] = 10'b0000000001;
assign label_8[849] = 10'b0000100000;
assign label_8[850] = 10'b0100000000;
assign label_8[851] = 10'b0010000000;
assign label_8[852] = 10'b1000000000;
assign label_8[853] = 10'b0000000100;
assign label_8[854] = 10'b0000010000;
assign label_8[855] = 10'b0001000000;
assign label_8[856] = 10'b0000000001;
assign label_8[857] = 10'b0000000001;
assign label_8[858] = 10'b0000010000;
assign label_8[859] = 10'b0000000001;
assign label_8[860] = 10'b0100000000;
assign label_8[861] = 10'b0100000000;
assign label_8[862] = 10'b1000000000;
assign label_8[863] = 10'b1000000000;
assign label_8[864] = 10'b0000100000;
assign label_8[865] = 10'b0000001000;
assign label_8[866] = 10'b0000000100;
assign label_8[867] = 10'b0001000000;
assign label_8[868] = 10'b0000000001;
assign label_8[869] = 10'b0001000000;
assign label_8[870] = 10'b0001000000;
assign label_8[871] = 10'b0000000001;
assign label_8[872] = 10'b0000100000;
assign label_8[873] = 10'b0000100000;
assign label_8[874] = 10'b0000100000;
assign label_8[875] = 10'b0000100000;
assign label_8[876] = 10'b0000100000;
assign label_8[877] = 10'b0100000000;
assign label_8[878] = 10'b0100000000;
assign label_8[879] = 10'b0100000000;
assign label_8[880] = 10'b0000100000;
assign label_8[881] = 10'b0000100000;
assign label_8[882] = 10'b0000010000;
assign label_8[883] = 10'b1000000000;
assign label_8[884] = 10'b0000010000;
assign label_8[885] = 10'b0000000001;
assign label_8[886] = 10'b0000000001;
assign label_8[887] = 10'b0000000001;
assign label_8[888] = 10'b0000000001;
assign label_8[889] = 10'b0000000001;
assign label_8[890] = 10'b0000010000;
assign label_8[891] = 10'b0000000100;
assign label_8[892] = 10'b0100000000;
assign label_8[893] = 10'b1000000000;
assign label_8[894] = 10'b0000000100;
assign label_8[895] = 10'b0000000100;
assign label_8[896] = 10'b0000000001;
assign label_8[897] = 10'b0000000100;
assign label_8[898] = 10'b0000100000;
assign label_8[899] = 10'b0000001000;
assign label_8[900] = 10'b0000001000;
assign label_8[901] = 10'b0000001000;
assign label_8[902] = 10'b0000000100;
assign label_8[903] = 10'b0000000100;
assign label_8[904] = 10'b0000000100;
assign label_8[905] = 10'b0000000100;
assign label_8[906] = 10'b0000000100;
assign label_8[907] = 10'b0000000100;
assign label_8[908] = 10'b0000000001;
assign label_8[909] = 10'b0100000000;
assign label_8[910] = 10'b0000001000;
assign label_8[911] = 10'b0000000100;
assign label_8[912] = 10'b0000000001;
assign label_8[913] = 10'b1000000000;
assign label_8[914] = 10'b0000000001;
assign label_8[915] = 10'b0000000100;
assign label_8[916] = 10'b0000100000;
assign label_8[917] = 10'b0000000001;
assign label_8[918] = 10'b0000000001;
assign label_8[919] = 10'b0000000001;
assign label_8[920] = 10'b0100000000;
assign label_8[921] = 10'b0000001000;
assign label_8[922] = 10'b0000000001;
assign label_8[923] = 10'b1000000000;
assign label_8[924] = 10'b0001000000;
assign label_8[925] = 10'b0001000000;
assign label_8[926] = 10'b0001000000;
assign label_8[927] = 10'b0001000000;
assign label_8[928] = 10'b0000010000;
assign label_8[929] = 10'b0000000001;
assign label_8[930] = 10'b0000100000;
assign label_8[931] = 10'b0001000000;
assign label_8[932] = 10'b0001000000;
assign label_8[933] = 10'b0000000001;
assign label_8[934] = 10'b0000000001;
assign label_8[935] = 10'b0001000000;
assign label_8[936] = 10'b0000000001;
assign label_8[937] = 10'b0000010000;
assign label_8[938] = 10'b1000000000;
assign label_8[939] = 10'b0000000001;
assign label_8[940] = 10'b0000000001;
assign label_8[941] = 10'b0000010000;
assign label_8[942] = 10'b0000000001;
assign label_8[943] = 10'b0000000001;
assign label_8[944] = 10'b0100000000;
assign label_8[945] = 10'b0000100000;
assign label_8[946] = 10'b0001000000;
assign label_8[947] = 10'b0100000000;
assign label_8[948] = 10'b0100000000;
assign label_8[949] = 10'b0100000000;
assign label_8[950] = 10'b0100000000;
assign label_8[951] = 10'b0000001000;
assign label_8[952] = 10'b0100000000;
assign label_8[953] = 10'b0000001000;
assign label_8[954] = 10'b0000000100;
assign label_8[955] = 10'b0000000100;
assign label_8[956] = 10'b0001000000;
assign label_8[957] = 10'b0000000001;
assign label_8[958] = 10'b0000000001;
assign label_8[959] = 10'b0000000001;
assign label_8[960] = 10'b0000010000;
assign label_8[961] = 10'b0010000000;
assign label_8[962] = 10'b0100000000;
assign label_8[963] = 10'b0001000000;
assign label_8[964] = 10'b0000100000;
assign label_8[965] = 10'b0001000000;
assign label_8[966] = 10'b0000000001;
assign label_8[967] = 10'b0000000001;
assign label_8[968] = 10'b0000010000;
assign label_8[969] = 10'b0000000100;
assign label_8[970] = 10'b0000010000;
assign label_8[971] = 10'b0001000000;
assign label_8[972] = 10'b0000000100;
assign label_8[973] = 10'b0000000100;
assign label_8[974] = 10'b0001000000;
assign label_8[975] = 10'b0001000000;
assign label_8[976] = 10'b0000000100;
assign label_8[977] = 10'b1000000000;
assign label_8[978] = 10'b1000000000;
assign label_8[979] = 10'b0000010000;
assign label_8[980] = 10'b0010000000;
assign label_8[981] = 10'b1000000000;
assign label_8[982] = 10'b0100000000;
assign label_8[983] = 10'b0100000000;
assign label_8[984] = 10'b0000010000;
assign label_8[985] = 10'b1000000000;
assign label_8[986] = 10'b0100000000;
assign label_8[987] = 10'b0000010000;
assign label_8[988] = 10'b0000010000;
assign label_8[989] = 10'b0000000100;
assign label_8[990] = 10'b0000000100;
assign label_8[991] = 10'b0000000100;
assign label_8[992] = 10'b0000000100;
assign label_8[993] = 10'b0010000000;
assign label_8[994] = 10'b0000000100;
assign label_8[995] = 10'b0001000000;
assign label_8[996] = 10'b0000000100;
assign label_8[997] = 10'b0000000100;
assign label_8[998] = 10'b0000000001;
assign label_8[999] = 10'b0001000000;
assign label_8[1000] = 10'b0000100000;
assign label_8[1001] = 10'b0100000000;
assign label_8[1002] = 10'b0000000100;
assign label_8[1003] = 10'b0000000100;
assign label_8[1004] = 10'b0100000000;
assign label_8[1005] = 10'b0100000000;
assign label_8[1006] = 10'b0001000000;
assign label_8[1007] = 10'b0001000000;
assign label_8[1008] = 10'b0000000100;
assign label_8[1009] = 10'b0000000100;
assign label_8[1010] = 10'b0000010000;
assign label_8[1011] = 10'b0100000000;
assign label_8[1012] = 10'b0000010000;
assign label_8[1013] = 10'b0100000000;
assign label_8[1014] = 10'b0100000000;
assign label_8[1015] = 10'b0001000000;
assign label_8[1016] = 10'b0000010000;
assign label_8[1017] = 10'b0000100000;
assign label_8[1018] = 10'b0000000001;
assign label_8[1019] = 10'b0000000100;
assign label_8[1020] = 10'b0000000001;
assign label_8[1021] = 10'b0100000000;
assign label_8[1022] = 10'b0001000000;
assign label_8[1023] = 10'b0000000001;
assign label_9[0] = 10'b1000000000;
assign label_9[1] = 10'b0000001000;
assign label_9[2] = 10'b0000000100;
assign label_9[3] = 10'b0001000000;
assign label_9[4] = 10'b0000100000;
assign label_9[5] = 10'b0000000001;
assign label_9[6] = 10'b0000100000;
assign label_9[7] = 10'b0000100000;
assign label_9[8] = 10'b0000000100;
assign label_9[9] = 10'b0000000100;
assign label_9[10] = 10'b0001000000;
assign label_9[11] = 10'b0000100000;
assign label_9[12] = 10'b0001000000;
assign label_9[13] = 10'b0001000000;
assign label_9[14] = 10'b0001000000;
assign label_9[15] = 10'b0000000010;
assign label_9[16] = 10'b0001000000;
assign label_9[17] = 10'b0001000000;
assign label_9[18] = 10'b0001000000;
assign label_9[19] = 10'b0000000100;
assign label_9[20] = 10'b0000000001;
assign label_9[21] = 10'b0000000001;
assign label_9[22] = 10'b0000010000;
assign label_9[23] = 10'b0000010000;
assign label_9[24] = 10'b0000000100;
assign label_9[25] = 10'b0000000100;
assign label_9[26] = 10'b0000000100;
assign label_9[27] = 10'b0001000000;
assign label_9[28] = 10'b0001000000;
assign label_9[29] = 10'b0001000000;
assign label_9[30] = 10'b0000000100;
assign label_9[31] = 10'b0001000000;
assign label_9[32] = 10'b0000010000;
assign label_9[33] = 10'b1000000000;
assign label_9[34] = 10'b0100000000;
assign label_9[35] = 10'b0000001000;
assign label_9[36] = 10'b1000000000;
assign label_9[37] = 10'b1000000000;
assign label_9[38] = 10'b0010000000;
assign label_9[39] = 10'b0000000100;
assign label_9[40] = 10'b0000010000;
assign label_9[41] = 10'b0001000000;
assign label_9[42] = 10'b0000010000;
assign label_9[43] = 10'b0000000100;
assign label_9[44] = 10'b0000000100;
assign label_9[45] = 10'b0000000100;
assign label_9[46] = 10'b0001000000;
assign label_9[47] = 10'b0000000100;
assign label_9[48] = 10'b0010000000;
assign label_9[49] = 10'b0010000000;
assign label_9[50] = 10'b0010000000;
assign label_9[51] = 10'b0000100000;
assign label_9[52] = 10'b0100000000;
assign label_9[53] = 10'b0000100000;
assign label_9[54] = 10'b0000000001;
assign label_9[55] = 10'b0000001000;
assign label_9[56] = 10'b0010000000;
assign label_9[57] = 10'b1000000000;
assign label_9[58] = 10'b1000000000;
assign label_9[59] = 10'b1000000000;
assign label_9[60] = 10'b0001000000;
assign label_9[61] = 10'b0000000001;
assign label_9[62] = 10'b0000000001;
assign label_9[63] = 10'b0000000100;
assign label_9[64] = 10'b0010000000;
assign label_9[65] = 10'b0010000000;
assign label_9[66] = 10'b0010000000;
assign label_9[67] = 10'b0010000000;
assign label_9[68] = 10'b1000000000;
assign label_9[69] = 10'b1000000000;
assign label_9[70] = 10'b1000000000;
assign label_9[71] = 10'b1000000000;
assign label_9[72] = 10'b0000100000;
assign label_9[73] = 10'b0000100000;
assign label_9[74] = 10'b0000100000;
assign label_9[75] = 10'b0000100000;
assign label_9[76] = 10'b1000000000;
assign label_9[77] = 10'b1000000000;
assign label_9[78] = 10'b1000000000;
assign label_9[79] = 10'b1000000000;
assign label_9[80] = 10'b0010000000;
assign label_9[81] = 10'b0010000000;
assign label_9[82] = 10'b0010000000;
assign label_9[83] = 10'b0010000000;
assign label_9[84] = 10'b0000010000;
assign label_9[85] = 10'b0000001000;
assign label_9[86] = 10'b0010000000;
assign label_9[87] = 10'b1000000000;
assign label_9[88] = 10'b0010000000;
assign label_9[89] = 10'b0010000000;
assign label_9[90] = 10'b1000000000;
assign label_9[91] = 10'b1000000000;
assign label_9[92] = 10'b1000000000;
assign label_9[93] = 10'b1000000000;
assign label_9[94] = 10'b0000010000;
assign label_9[95] = 10'b1000000000;
assign label_9[96] = 10'b1000000000;
assign label_9[97] = 10'b0010000000;
assign label_9[98] = 10'b0010000000;
assign label_9[99] = 10'b0010000000;
assign label_9[100] = 10'b1000000000;
assign label_9[101] = 10'b1000000000;
assign label_9[102] = 10'b0000100000;
assign label_9[103] = 10'b1000000000;
assign label_9[104] = 10'b0000010000;
assign label_9[105] = 10'b0000010000;
assign label_9[106] = 10'b0000010000;
assign label_9[107] = 10'b0000010000;
assign label_9[108] = 10'b0010000000;
assign label_9[109] = 10'b0010000000;
assign label_9[110] = 10'b0010000000;
assign label_9[111] = 10'b0010000000;
assign label_9[112] = 10'b0010000000;
assign label_9[113] = 10'b0010000000;
assign label_9[114] = 10'b0010000000;
assign label_9[115] = 10'b0010000000;
assign label_9[116] = 10'b0010000000;
assign label_9[117] = 10'b0010000000;
assign label_9[118] = 10'b0010000000;
assign label_9[119] = 10'b0010000000;
assign label_9[120] = 10'b1000000000;
assign label_9[121] = 10'b1000000000;
assign label_9[122] = 10'b1000000000;
assign label_9[123] = 10'b1000000000;
assign label_9[124] = 10'b1000000000;
assign label_9[125] = 10'b1000000000;
assign label_9[126] = 10'b1000000000;
assign label_9[127] = 10'b1000000000;
assign label_9[128] = 10'b0000000001;
assign label_9[129] = 10'b0010000000;
assign label_9[130] = 10'b0000000001;
assign label_9[131] = 10'b0000000100;
assign label_9[132] = 10'b0001000000;
assign label_9[133] = 10'b0000100000;
assign label_9[134] = 10'b0000100000;
assign label_9[135] = 10'b0100000000;
assign label_9[136] = 10'b0001000000;
assign label_9[137] = 10'b0010000000;
assign label_9[138] = 10'b1000000000;
assign label_9[139] = 10'b0000000001;
assign label_9[140] = 10'b0000000100;
assign label_9[141] = 10'b0000001000;
assign label_9[142] = 10'b0000000100;
assign label_9[143] = 10'b0000000001;
assign label_9[144] = 10'b0000001000;
assign label_9[145] = 10'b0000100000;
assign label_9[146] = 10'b0100000000;
assign label_9[147] = 10'b0001000000;
assign label_9[148] = 10'b0000001000;
assign label_9[149] = 10'b1000000000;
assign label_9[150] = 10'b0000000100;
assign label_9[151] = 10'b0100000000;
assign label_9[152] = 10'b0000100000;
assign label_9[153] = 10'b0000100000;
assign label_9[154] = 10'b0000100000;
assign label_9[155] = 10'b0000100000;
assign label_9[156] = 10'b0000100000;
assign label_9[157] = 10'b0000001000;
assign label_9[158] = 10'b0100000000;
assign label_9[159] = 10'b0000100000;
assign label_9[160] = 10'b0000001000;
assign label_9[161] = 10'b0000100000;
assign label_9[162] = 10'b0001000000;
assign label_9[163] = 10'b0100000000;
assign label_9[164] = 10'b0000100000;
assign label_9[165] = 10'b0001000000;
assign label_9[166] = 10'b0000001000;
assign label_9[167] = 10'b0000100000;
assign label_9[168] = 10'b0000001000;
assign label_9[169] = 10'b0000100000;
assign label_9[170] = 10'b0000001000;
assign label_9[171] = 10'b0000100000;
assign label_9[172] = 10'b0001000000;
assign label_9[173] = 10'b0000000001;
assign label_9[174] = 10'b0010000000;
assign label_9[175] = 10'b0000000001;
assign label_9[176] = 10'b0000001000;
assign label_9[177] = 10'b0010000000;
assign label_9[178] = 10'b0000001000;
assign label_9[179] = 10'b0000001000;
assign label_9[180] = 10'b0000001000;
assign label_9[181] = 10'b0000001000;
assign label_9[182] = 10'b0000000100;
assign label_9[183] = 10'b0000001000;
assign label_9[184] = 10'b0100000000;
assign label_9[185] = 10'b0000000100;
assign label_9[186] = 10'b0000000100;
assign label_9[187] = 10'b0000001000;
assign label_9[188] = 10'b0000000100;
assign label_9[189] = 10'b0000000100;
assign label_9[190] = 10'b0100000000;
assign label_9[191] = 10'b0000001000;
assign label_9[192] = 10'b0000000001;
assign label_9[193] = 10'b0000100000;
assign label_9[194] = 10'b0000000001;
assign label_9[195] = 10'b0000000001;
assign label_9[196] = 10'b0000100000;
assign label_9[197] = 10'b0100000000;
assign label_9[198] = 10'b0010000000;
assign label_9[199] = 10'b1000000000;
assign label_9[200] = 10'b0000100000;
assign label_9[201] = 10'b0000100000;
assign label_9[202] = 10'b0000100000;
assign label_9[203] = 10'b0000001000;
assign label_9[204] = 10'b0000100000;
assign label_9[205] = 10'b0100000000;
assign label_9[206] = 10'b0001000000;
assign label_9[207] = 10'b0000001000;
assign label_9[208] = 10'b0000000001;
assign label_9[209] = 10'b0000000001;
assign label_9[210] = 10'b0000000001;
assign label_9[211] = 10'b0000000001;
assign label_9[212] = 10'b0000000001;
assign label_9[213] = 10'b0000000001;
assign label_9[214] = 10'b0001000000;
assign label_9[215] = 10'b0001000000;
assign label_9[216] = 10'b0000000001;
assign label_9[217] = 10'b0000000001;
assign label_9[218] = 10'b0000000001;
assign label_9[219] = 10'b0000000001;
assign label_9[220] = 10'b0000100000;
assign label_9[221] = 10'b0000100000;
assign label_9[222] = 10'b0000100000;
assign label_9[223] = 10'b0000100000;
assign label_9[224] = 10'b0010000000;
assign label_9[225] = 10'b0010000000;
assign label_9[226] = 10'b1000000000;
assign label_9[227] = 10'b1000000000;
assign label_9[228] = 10'b1000000000;
assign label_9[229] = 10'b1000000000;
assign label_9[230] = 10'b0000001000;
assign label_9[231] = 10'b0000001000;
assign label_9[232] = 10'b0010000000;
assign label_9[233] = 10'b0010000000;
assign label_9[234] = 10'b1000000000;
assign label_9[235] = 10'b0010000000;
assign label_9[236] = 10'b1000000000;
assign label_9[237] = 10'b1000000000;
assign label_9[238] = 10'b0000100000;
assign label_9[239] = 10'b0000100000;
assign label_9[240] = 10'b0000100000;
assign label_9[241] = 10'b0000100000;
assign label_9[242] = 10'b0000001000;
assign label_9[243] = 10'b0000100000;
assign label_9[244] = 10'b1000000000;
assign label_9[245] = 10'b0000001000;
assign label_9[246] = 10'b0000100000;
assign label_9[247] = 10'b0000001000;
assign label_9[248] = 10'b0000001000;
assign label_9[249] = 10'b0000001000;
assign label_9[250] = 10'b1000000000;
assign label_9[251] = 10'b1000000000;
assign label_9[252] = 10'b1000000000;
assign label_9[253] = 10'b0010000000;
assign label_9[254] = 10'b1000000000;
assign label_9[255] = 10'b0010000000;
assign label_9[256] = 10'b0000100000;
assign label_9[257] = 10'b0010000000;
assign label_9[258] = 10'b0001000000;
assign label_9[259] = 10'b0010000000;
assign label_9[260] = 10'b0000000001;
assign label_9[261] = 10'b0000000001;
assign label_9[262] = 10'b0010000000;
assign label_9[263] = 10'b0010000000;
assign label_9[264] = 10'b0010000000;
assign label_9[265] = 10'b0001000000;
assign label_9[266] = 10'b1000000000;
assign label_9[267] = 10'b0000001000;
assign label_9[268] = 10'b0000100000;
assign label_9[269] = 10'b0100000000;
assign label_9[270] = 10'b0000100000;
assign label_9[271] = 10'b1000000000;
assign label_9[272] = 10'b0100000000;
assign label_9[273] = 10'b0000010000;
assign label_9[274] = 10'b0001000000;
assign label_9[275] = 10'b0001000000;
assign label_9[276] = 10'b0010000000;
assign label_9[277] = 10'b0010000000;
assign label_9[278] = 10'b0010000000;
assign label_9[279] = 10'b0010000000;
assign label_9[280] = 10'b0000000001;
assign label_9[281] = 10'b0000001000;
assign label_9[282] = 10'b0000000100;
assign label_9[283] = 10'b0000100000;
assign label_9[284] = 10'b0000001000;
assign label_9[285] = 10'b0000001000;
assign label_9[286] = 10'b0100000000;
assign label_9[287] = 10'b0100000000;
assign label_9[288] = 10'b0010000000;
assign label_9[289] = 10'b0010000000;
assign label_9[290] = 10'b0000000001;
assign label_9[291] = 10'b0000000100;
assign label_9[292] = 10'b0000010000;
assign label_9[293] = 10'b1000000000;
assign label_9[294] = 10'b0000100000;
assign label_9[295] = 10'b0000010000;
assign label_9[296] = 10'b0000000001;
assign label_9[297] = 10'b0000000001;
assign label_9[298] = 10'b0000001000;
assign label_9[299] = 10'b0000000100;
assign label_9[300] = 10'b0000000001;
assign label_9[301] = 10'b0000000001;
assign label_9[302] = 10'b0000001000;
assign label_9[303] = 10'b0000001000;
assign label_9[304] = 10'b1000000000;
assign label_9[305] = 10'b1000000000;
assign label_9[306] = 10'b0000010000;
assign label_9[307] = 10'b1000000000;
assign label_9[308] = 10'b0000001000;
assign label_9[309] = 10'b0000001000;
assign label_9[310] = 10'b0100000000;
assign label_9[311] = 10'b0100000000;
assign label_9[312] = 10'b0000010000;
assign label_9[313] = 10'b1000000000;
assign label_9[314] = 10'b0000100000;
assign label_9[315] = 10'b0000001000;
assign label_9[316] = 10'b0000001000;
assign label_9[317] = 10'b0000100000;
assign label_9[318] = 10'b0000001000;
assign label_9[319] = 10'b1000000000;
assign label_9[320] = 10'b0000000001;
assign label_9[321] = 10'b0000000100;
assign label_9[322] = 10'b0000000001;
assign label_9[323] = 10'b0000000001;
assign label_9[324] = 10'b0000000001;
assign label_9[325] = 10'b0000000001;
assign label_9[326] = 10'b0000000100;
assign label_9[327] = 10'b0000100000;
assign label_9[328] = 10'b0100000000;
assign label_9[329] = 10'b0100000000;
assign label_9[330] = 10'b0000100000;
assign label_9[331] = 10'b0000100000;
assign label_9[332] = 10'b0000000001;
assign label_9[333] = 10'b0000000001;
assign label_9[334] = 10'b0000000001;
assign label_9[335] = 10'b0000000001;
assign label_9[336] = 10'b0000000001;
assign label_9[337] = 10'b0000000100;
assign label_9[338] = 10'b0000000100;
assign label_9[339] = 10'b0000000001;
assign label_9[340] = 10'b0000001000;
assign label_9[341] = 10'b0000001000;
assign label_9[342] = 10'b0000000001;
assign label_9[343] = 10'b0000100000;
assign label_9[344] = 10'b0000000100;
assign label_9[345] = 10'b0000000100;
assign label_9[346] = 10'b0000000100;
assign label_9[347] = 10'b0000000100;
assign label_9[348] = 10'b0000000001;
assign label_9[349] = 10'b0000000001;
assign label_9[350] = 10'b0000000001;
assign label_9[351] = 10'b0000000100;
assign label_9[352] = 10'b0000001000;
assign label_9[353] = 10'b0100000000;
assign label_9[354] = 10'b0000001000;
assign label_9[355] = 10'b0000001000;
assign label_9[356] = 10'b0000010000;
assign label_9[357] = 10'b0000100000;
assign label_9[358] = 10'b0100000000;
assign label_9[359] = 10'b0000001000;
assign label_9[360] = 10'b0000001000;
assign label_9[361] = 10'b0000100000;
assign label_9[362] = 10'b0000001000;
assign label_9[363] = 10'b0000001000;
assign label_9[364] = 10'b0000001000;
assign label_9[365] = 10'b0000100000;
assign label_9[366] = 10'b0000001000;
assign label_9[367] = 10'b1000000000;
assign label_9[368] = 10'b0100000000;
assign label_9[369] = 10'b0000000100;
assign label_9[370] = 10'b0100000000;
assign label_9[371] = 10'b0100000000;
assign label_9[372] = 10'b0100000000;
assign label_9[373] = 10'b0100000000;
assign label_9[374] = 10'b0100000000;
assign label_9[375] = 10'b0100000000;
assign label_9[376] = 10'b0000000001;
assign label_9[377] = 10'b1000000000;
assign label_9[378] = 10'b0100000000;
assign label_9[379] = 10'b0000000100;
assign label_9[380] = 10'b0000000001;
assign label_9[381] = 10'b0100000000;
assign label_9[382] = 10'b0000001000;
assign label_9[383] = 10'b0000001000;
assign label_9[384] = 10'b0010000000;
assign label_9[385] = 10'b0000000001;
assign label_9[386] = 10'b0000010000;
assign label_9[387] = 10'b0000010000;
assign label_9[388] = 10'b0000100000;
assign label_9[389] = 10'b0000010000;
assign label_9[390] = 10'b0001000000;
assign label_9[391] = 10'b0000000001;
assign label_9[392] = 10'b1000000000;
assign label_9[393] = 10'b0010000000;
assign label_9[394] = 10'b0000000001;
assign label_9[395] = 10'b0010000000;
assign label_9[396] = 10'b0000001000;
assign label_9[397] = 10'b1000000000;
assign label_9[398] = 10'b0000001000;
assign label_9[399] = 10'b1000000000;
assign label_9[400] = 10'b0000100000;
assign label_9[401] = 10'b0000010000;
assign label_9[402] = 10'b0000000001;
assign label_9[403] = 10'b0000000100;
assign label_9[404] = 10'b0000000001;
assign label_9[405] = 10'b0000000001;
assign label_9[406] = 10'b0010000000;
assign label_9[407] = 10'b0010000000;
assign label_9[408] = 10'b0000010000;
assign label_9[409] = 10'b0000010000;
assign label_9[410] = 10'b0000010000;
assign label_9[411] = 10'b0000010000;
assign label_9[412] = 10'b0010000000;
assign label_9[413] = 10'b0010000000;
assign label_9[414] = 10'b0010000000;
assign label_9[415] = 10'b0010000000;
assign label_9[416] = 10'b1000000000;
assign label_9[417] = 10'b1000000000;
assign label_9[418] = 10'b1000000000;
assign label_9[419] = 10'b1000000000;
assign label_9[420] = 10'b0000010000;
assign label_9[421] = 10'b0000000100;
assign label_9[422] = 10'b1000000000;
assign label_9[423] = 10'b0000000001;
assign label_9[424] = 10'b0000000100;
assign label_9[425] = 10'b0000000100;
assign label_9[426] = 10'b0000010000;
assign label_9[427] = 10'b0000010000;
assign label_9[428] = 10'b0000000001;
assign label_9[429] = 10'b1000000000;
assign label_9[430] = 10'b0001000000;
assign label_9[431] = 10'b0001000000;
assign label_9[432] = 10'b0000000001;
assign label_9[433] = 10'b0000000001;
assign label_9[434] = 10'b0000000001;
assign label_9[435] = 10'b0100000000;
assign label_9[436] = 10'b0100000000;
assign label_9[437] = 10'b0000001000;
assign label_9[438] = 10'b0000000001;
assign label_9[439] = 10'b0100000000;
assign label_9[440] = 10'b0000010000;
assign label_9[441] = 10'b0000010000;
assign label_9[442] = 10'b0000010000;
assign label_9[443] = 10'b0000010000;
assign label_9[444] = 10'b0010000000;
assign label_9[445] = 10'b0010000000;
assign label_9[446] = 10'b1000000000;
assign label_9[447] = 10'b1000000000;
assign label_9[448] = 10'b0000000001;
assign label_9[449] = 10'b0000000001;
assign label_9[450] = 10'b0000000100;
assign label_9[451] = 10'b0000000100;
assign label_9[452] = 10'b0000000001;
assign label_9[453] = 10'b0000000001;
assign label_9[454] = 10'b1000000000;
assign label_9[455] = 10'b0000100000;
assign label_9[456] = 10'b0000100000;
assign label_9[457] = 10'b0100000000;
assign label_9[458] = 10'b0001000000;
assign label_9[459] = 10'b0000000001;
assign label_9[460] = 10'b0000000100;
assign label_9[461] = 10'b0000000100;
assign label_9[462] = 10'b0000000001;
assign label_9[463] = 10'b0001000000;
assign label_9[464] = 10'b0000010000;
assign label_9[465] = 10'b0000000100;
assign label_9[466] = 10'b0100000000;
assign label_9[467] = 10'b0001000000;
assign label_9[468] = 10'b0001000000;
assign label_9[469] = 10'b0001000000;
assign label_9[470] = 10'b0000000100;
assign label_9[471] = 10'b0001000000;
assign label_9[472] = 10'b0000100000;
assign label_9[473] = 10'b0000100000;
assign label_9[474] = 10'b0000000001;
assign label_9[475] = 10'b0000000001;
assign label_9[476] = 10'b0010000000;
assign label_9[477] = 10'b0000000001;
assign label_9[478] = 10'b0000000001;
assign label_9[479] = 10'b0000000001;
assign label_9[480] = 10'b0000000001;
assign label_9[481] = 10'b0000000001;
assign label_9[482] = 10'b0000000100;
assign label_9[483] = 10'b0000000001;
assign label_9[484] = 10'b0000000100;
assign label_9[485] = 10'b0100000000;
assign label_9[486] = 10'b0000000001;
assign label_9[487] = 10'b0000001000;
assign label_9[488] = 10'b0000000001;
assign label_9[489] = 10'b0000000001;
assign label_9[490] = 10'b0000000001;
assign label_9[491] = 10'b0000000001;
assign label_9[492] = 10'b0000000100;
assign label_9[493] = 10'b0000000100;
assign label_9[494] = 10'b0000000100;
assign label_9[495] = 10'b0000000100;
assign label_9[496] = 10'b1000000000;
assign label_9[497] = 10'b1000000000;
assign label_9[498] = 10'b1000000000;
assign label_9[499] = 10'b1000000000;
assign label_9[500] = 10'b0000001000;
assign label_9[501] = 10'b0000000100;
assign label_9[502] = 10'b0000000001;
assign label_9[503] = 10'b0100000000;
assign label_9[504] = 10'b0100000000;
assign label_9[505] = 10'b0000000001;
assign label_9[506] = 10'b0000001000;
assign label_9[507] = 10'b0000000100;
assign label_9[508] = 10'b0001000000;
assign label_9[509] = 10'b0000000001;
assign label_9[510] = 10'b1000000000;
assign label_9[511] = 10'b0000000001;
assign label_9[512] = 10'b0000000010;
assign label_9[513] = 10'b0000010000;
assign label_9[514] = 10'b0000001000;
assign label_9[515] = 10'b0000000010;
assign label_9[516] = 10'b0010000000;
assign label_9[517] = 10'b0100000000;
assign label_9[518] = 10'b1000000000;
assign label_9[519] = 10'b0100000000;
assign label_9[520] = 10'b0000000100;
assign label_9[521] = 10'b0000001000;
assign label_9[522] = 10'b0000000100;
assign label_9[523] = 10'b0000100000;
assign label_9[524] = 10'b0010000000;
assign label_9[525] = 10'b0000001000;
assign label_9[526] = 10'b0010000000;
assign label_9[527] = 10'b0000001000;
assign label_9[528] = 10'b0000001000;
assign label_9[529] = 10'b0000001000;
assign label_9[530] = 10'b1000000000;
assign label_9[531] = 10'b0000010000;
assign label_9[532] = 10'b0000010000;
assign label_9[533] = 10'b0010000000;
assign label_9[534] = 10'b0100000000;
assign label_9[535] = 10'b0000000100;
assign label_9[536] = 10'b0001000000;
assign label_9[537] = 10'b0000000100;
assign label_9[538] = 10'b0000000100;
assign label_9[539] = 10'b0100000000;
assign label_9[540] = 10'b0001000000;
assign label_9[541] = 10'b0000000100;
assign label_9[542] = 10'b0010000000;
assign label_9[543] = 10'b0000000010;
assign label_9[544] = 10'b0010000000;
assign label_9[545] = 10'b0000000100;
assign label_9[546] = 10'b0000100000;
assign label_9[547] = 10'b0000000100;
assign label_9[548] = 10'b0010000000;
assign label_9[549] = 10'b0000000100;
assign label_9[550] = 10'b0010000000;
assign label_9[551] = 10'b0000000100;
assign label_9[552] = 10'b0010000000;
assign label_9[553] = 10'b0000010000;
assign label_9[554] = 10'b0000010000;
assign label_9[555] = 10'b0000100000;
assign label_9[556] = 10'b0000000100;
assign label_9[557] = 10'b0000000100;
assign label_9[558] = 10'b0000100000;
assign label_9[559] = 10'b0000100000;
assign label_9[560] = 10'b0010000000;
assign label_9[561] = 10'b0000001000;
assign label_9[562] = 10'b0000001000;
assign label_9[563] = 10'b0000001000;
assign label_9[564] = 10'b0100000000;
assign label_9[565] = 10'b0100000000;
assign label_9[566] = 10'b0000000010;
assign label_9[567] = 10'b0010000000;
assign label_9[568] = 10'b0010000000;
assign label_9[569] = 10'b0100000000;
assign label_9[570] = 10'b0000100000;
assign label_9[571] = 10'b0100000000;
assign label_9[572] = 10'b0000100000;
assign label_9[573] = 10'b0000100000;
assign label_9[574] = 10'b0100000000;
assign label_9[575] = 10'b0100000000;
assign label_9[576] = 10'b0000010000;
assign label_9[577] = 10'b1000000000;
assign label_9[578] = 10'b1000000000;
assign label_9[579] = 10'b1000000000;
assign label_9[580] = 10'b0000000100;
assign label_9[581] = 10'b0010000000;
assign label_9[582] = 10'b0001000000;
assign label_9[583] = 10'b0000010000;
assign label_9[584] = 10'b0000100000;
assign label_9[585] = 10'b0100000000;
assign label_9[586] = 10'b0000010000;
assign label_9[587] = 10'b0001000000;
assign label_9[588] = 10'b0001000000;
assign label_9[589] = 10'b0001000000;
assign label_9[590] = 10'b0001000000;
assign label_9[591] = 10'b0001000000;
assign label_9[592] = 10'b0010000000;
assign label_9[593] = 10'b1000000000;
assign label_9[594] = 10'b1000000000;
assign label_9[595] = 10'b0100000000;
assign label_9[596] = 10'b0010000000;
assign label_9[597] = 10'b0000001000;
assign label_9[598] = 10'b0000001000;
assign label_9[599] = 10'b0100000000;
assign label_9[600] = 10'b0010000000;
assign label_9[601] = 10'b0000100000;
assign label_9[602] = 10'b0000100000;
assign label_9[603] = 10'b0010000000;
assign label_9[604] = 10'b0100000000;
assign label_9[605] = 10'b0100000000;
assign label_9[606] = 10'b0010000000;
assign label_9[607] = 10'b0010000000;
assign label_9[608] = 10'b0000100000;
assign label_9[609] = 10'b0000100000;
assign label_9[610] = 10'b0000100000;
assign label_9[611] = 10'b0100000000;
assign label_9[612] = 10'b1000000000;
assign label_9[613] = 10'b0100000000;
assign label_9[614] = 10'b0100000000;
assign label_9[615] = 10'b0001000000;
assign label_9[616] = 10'b0100000000;
assign label_9[617] = 10'b0000100000;
assign label_9[618] = 10'b1000000000;
assign label_9[619] = 10'b0000000010;
assign label_9[620] = 10'b0001000000;
assign label_9[621] = 10'b0100000000;
assign label_9[622] = 10'b0100000000;
assign label_9[623] = 10'b0100000000;
assign label_9[624] = 10'b1000000000;
assign label_9[625] = 10'b0010000000;
assign label_9[626] = 10'b1000000000;
assign label_9[627] = 10'b0100000000;
assign label_9[628] = 10'b0000010000;
assign label_9[629] = 10'b0100000000;
assign label_9[630] = 10'b0001000000;
assign label_9[631] = 10'b0100000000;
assign label_9[632] = 10'b0100000000;
assign label_9[633] = 10'b0000010000;
assign label_9[634] = 10'b0100000000;
assign label_9[635] = 10'b1000000000;
assign label_9[636] = 10'b0000010000;
assign label_9[637] = 10'b0100000000;
assign label_9[638] = 10'b0100000000;
assign label_9[639] = 10'b0100000000;
assign label_9[640] = 10'b0000010000;
assign label_9[641] = 10'b0001000000;
assign label_9[642] = 10'b0000010000;
assign label_9[643] = 10'b0000000100;
assign label_9[644] = 10'b0000100000;
assign label_9[645] = 10'b0000010000;
assign label_9[646] = 10'b0000010000;
assign label_9[647] = 10'b0000010000;
assign label_9[648] = 10'b0001000000;
assign label_9[649] = 10'b0001000000;
assign label_9[650] = 10'b0001000000;
assign label_9[651] = 10'b0001000000;
assign label_9[652] = 10'b0001000000;
assign label_9[653] = 10'b0001000000;
assign label_9[654] = 10'b0001000000;
assign label_9[655] = 10'b0001000000;
assign label_9[656] = 10'b0001000000;
assign label_9[657] = 10'b0001000000;
assign label_9[658] = 10'b0000010000;
assign label_9[659] = 10'b0001000000;
assign label_9[660] = 10'b0000000100;
assign label_9[661] = 10'b0000000100;
assign label_9[662] = 10'b0000000100;
assign label_9[663] = 10'b0000000100;
assign label_9[664] = 10'b0000000100;
assign label_9[665] = 10'b0000000100;
assign label_9[666] = 10'b0000000100;
assign label_9[667] = 10'b0000000100;
assign label_9[668] = 10'b0000000100;
assign label_9[669] = 10'b0000000100;
assign label_9[670] = 10'b0000000100;
assign label_9[671] = 10'b0000000100;
assign label_9[672] = 10'b0010000000;
assign label_9[673] = 10'b0010000000;
assign label_9[674] = 10'b0000010000;
assign label_9[675] = 10'b0000010000;
assign label_9[676] = 10'b1000000000;
assign label_9[677] = 10'b0000010000;
assign label_9[678] = 10'b0000010000;
assign label_9[679] = 10'b0000010000;
assign label_9[680] = 10'b0010000000;
assign label_9[681] = 10'b0010000000;
assign label_9[682] = 10'b0010000000;
assign label_9[683] = 10'b0000010000;
assign label_9[684] = 10'b0000100000;
assign label_9[685] = 10'b1000000000;
assign label_9[686] = 10'b0010000000;
assign label_9[687] = 10'b0010000000;
assign label_9[688] = 10'b1000000000;
assign label_9[689] = 10'b0010000000;
assign label_9[690] = 10'b0010000000;
assign label_9[691] = 10'b0010000000;
assign label_9[692] = 10'b1000000000;
assign label_9[693] = 10'b0000010000;
assign label_9[694] = 10'b0000100000;
assign label_9[695] = 10'b0000100000;
assign label_9[696] = 10'b0000010000;
assign label_9[697] = 10'b0000010000;
assign label_9[698] = 10'b0000010000;
assign label_9[699] = 10'b0000010000;
assign label_9[700] = 10'b0000100000;
assign label_9[701] = 10'b0000100000;
assign label_9[702] = 10'b0010000000;
assign label_9[703] = 10'b0010000000;
assign label_9[704] = 10'b0000100000;
assign label_9[705] = 10'b1000000000;
assign label_9[706] = 10'b0000100000;
assign label_9[707] = 10'b0000000100;
assign label_9[708] = 10'b0000000100;
assign label_9[709] = 10'b0000000100;
assign label_9[710] = 10'b0000000100;
assign label_9[711] = 10'b0000000100;
assign label_9[712] = 10'b1000000000;
assign label_9[713] = 10'b0010000000;
assign label_9[714] = 10'b0000000100;
assign label_9[715] = 10'b0010000000;
assign label_9[716] = 10'b0000000100;
assign label_9[717] = 10'b0000010000;
assign label_9[718] = 10'b0001000000;
assign label_9[719] = 10'b0000010000;
assign label_9[720] = 10'b0000001000;
assign label_9[721] = 10'b0000000100;
assign label_9[722] = 10'b1000000000;
assign label_9[723] = 10'b0100000000;
assign label_9[724] = 10'b1000000000;
assign label_9[725] = 10'b0001000000;
assign label_9[726] = 10'b0100000000;
assign label_9[727] = 10'b0000100000;
assign label_9[728] = 10'b0000001000;
assign label_9[729] = 10'b0100000000;
assign label_9[730] = 10'b1000000000;
assign label_9[731] = 10'b0000010000;
assign label_9[732] = 10'b0000100000;
assign label_9[733] = 10'b0000001000;
assign label_9[734] = 10'b0000001000;
assign label_9[735] = 10'b0000001000;
assign label_9[736] = 10'b0000010000;
assign label_9[737] = 10'b0001000000;
assign label_9[738] = 10'b0000010000;
assign label_9[739] = 10'b0000100000;
assign label_9[740] = 10'b0000010000;
assign label_9[741] = 10'b0100000000;
assign label_9[742] = 10'b1000000000;
assign label_9[743] = 10'b0000010000;
assign label_9[744] = 10'b0000010000;
assign label_9[745] = 10'b0001000000;
assign label_9[746] = 10'b0001000000;
assign label_9[747] = 10'b0001000000;
assign label_9[748] = 10'b0000100000;
assign label_9[749] = 10'b0000010000;
assign label_9[750] = 10'b1000000000;
assign label_9[751] = 10'b1000000000;
assign label_9[752] = 10'b1000000000;
assign label_9[753] = 10'b1000000000;
assign label_9[754] = 10'b1000000000;
assign label_9[755] = 10'b0000100000;
assign label_9[756] = 10'b0000100000;
assign label_9[757] = 10'b0000100000;
assign label_9[758] = 10'b0000100000;
assign label_9[759] = 10'b0000100000;
assign label_9[760] = 10'b0000010000;
assign label_9[761] = 10'b0010000000;
assign label_9[762] = 10'b1000000000;
assign label_9[763] = 10'b0000010000;
assign label_9[764] = 10'b0000001000;
assign label_9[765] = 10'b0000001000;
assign label_9[766] = 10'b0010000000;
assign label_9[767] = 10'b0000100000;
assign label_9[768] = 10'b0010000000;
assign label_9[769] = 10'b0000000100;
assign label_9[770] = 10'b0000100000;
assign label_9[771] = 10'b0001000000;
assign label_9[772] = 10'b0000000010;
assign label_9[773] = 10'b0000000010;
assign label_9[774] = 10'b0000000010;
assign label_9[775] = 10'b0100000000;
assign label_9[776] = 10'b0000000100;
assign label_9[777] = 10'b0000010000;
assign label_9[778] = 10'b0001000000;
assign label_9[779] = 10'b0100000000;
assign label_9[780] = 10'b0001000000;
assign label_9[781] = 10'b0001000000;
assign label_9[782] = 10'b0001000000;
assign label_9[783] = 10'b0001000000;
assign label_9[784] = 10'b0001000000;
assign label_9[785] = 10'b0000000100;
assign label_9[786] = 10'b0001000000;
assign label_9[787] = 10'b0000001000;
assign label_9[788] = 10'b0010000000;
assign label_9[789] = 10'b0000100000;
assign label_9[790] = 10'b0100000000;
assign label_9[791] = 10'b0000100000;
assign label_9[792] = 10'b0001000000;
assign label_9[793] = 10'b0100000000;
assign label_9[794] = 10'b0000000100;
assign label_9[795] = 10'b0000010000;
assign label_9[796] = 10'b0000000100;
assign label_9[797] = 10'b0001000000;
assign label_9[798] = 10'b0001000000;
assign label_9[799] = 10'b0001000000;
assign label_9[800] = 10'b0000100000;
assign label_9[801] = 10'b0000100000;
assign label_9[802] = 10'b0000100000;
assign label_9[803] = 10'b0000100000;
assign label_9[804] = 10'b0000100000;
assign label_9[805] = 10'b0000001000;
assign label_9[806] = 10'b0000100000;
assign label_9[807] = 10'b0000100000;
assign label_9[808] = 10'b0000000001;
assign label_9[809] = 10'b0000001000;
assign label_9[810] = 10'b0100000000;
assign label_9[811] = 10'b0000100000;
assign label_9[812] = 10'b0100000000;
assign label_9[813] = 10'b0100000000;
assign label_9[814] = 10'b0100000000;
assign label_9[815] = 10'b0100000000;
assign label_9[816] = 10'b0000010000;
assign label_9[817] = 10'b0000100000;
assign label_9[818] = 10'b0001000000;
assign label_9[819] = 10'b0001000000;
assign label_9[820] = 10'b0000000100;
assign label_9[821] = 10'b0100000000;
assign label_9[822] = 10'b0000010000;
assign label_9[823] = 10'b0000010000;
assign label_9[824] = 10'b0000100000;
assign label_9[825] = 10'b0000100000;
assign label_9[826] = 10'b0100000000;
assign label_9[827] = 10'b0010000000;
assign label_9[828] = 10'b0010000000;
assign label_9[829] = 10'b0000010000;
assign label_9[830] = 10'b0100000000;
assign label_9[831] = 10'b0100000000;
assign label_9[832] = 10'b0000000100;
assign label_9[833] = 10'b0000000100;
assign label_9[834] = 10'b0000000100;
assign label_9[835] = 10'b0100000000;
assign label_9[836] = 10'b0001000000;
assign label_9[837] = 10'b0000000100;
assign label_9[838] = 10'b1000000000;
assign label_9[839] = 10'b1000000000;
assign label_9[840] = 10'b0100000000;
assign label_9[841] = 10'b0000000100;
assign label_9[842] = 10'b0010000000;
assign label_9[843] = 10'b1000000000;
assign label_9[844] = 10'b0000000100;
assign label_9[845] = 10'b0000000100;
assign label_9[846] = 10'b0100000000;
assign label_9[847] = 10'b0000000100;
assign label_9[848] = 10'b0100000000;
assign label_9[849] = 10'b0000000100;
assign label_9[850] = 10'b0100000000;
assign label_9[851] = 10'b0100000000;
assign label_9[852] = 10'b0000001000;
assign label_9[853] = 10'b0100000000;
assign label_9[854] = 10'b0000100000;
assign label_9[855] = 10'b0100000000;
assign label_9[856] = 10'b0000001000;
assign label_9[857] = 10'b0000000100;
assign label_9[858] = 10'b0000000100;
assign label_9[859] = 10'b0100000000;
assign label_9[860] = 10'b0000001000;
assign label_9[861] = 10'b0100000000;
assign label_9[862] = 10'b0000000100;
assign label_9[863] = 10'b0100000000;
assign label_9[864] = 10'b0001000000;
assign label_9[865] = 10'b0100000000;
assign label_9[866] = 10'b0000100000;
assign label_9[867] = 10'b0100000000;
assign label_9[868] = 10'b0000100000;
assign label_9[869] = 10'b0100000000;
assign label_9[870] = 10'b0000100000;
assign label_9[871] = 10'b0100000000;
assign label_9[872] = 10'b0001000000;
assign label_9[873] = 10'b0000000001;
assign label_9[874] = 10'b0100000000;
assign label_9[875] = 10'b0000000100;
assign label_9[876] = 10'b0000100000;
assign label_9[877] = 10'b0100000000;
assign label_9[878] = 10'b0100000000;
assign label_9[879] = 10'b0001000000;
assign label_9[880] = 10'b0000000100;
assign label_9[881] = 10'b1000000000;
assign label_9[882] = 10'b0100000000;
assign label_9[883] = 10'b0001000000;
assign label_9[884] = 10'b0001000000;
assign label_9[885] = 10'b0001000000;
assign label_9[886] = 10'b0001000000;
assign label_9[887] = 10'b0001000000;
assign label_9[888] = 10'b0100000000;
assign label_9[889] = 10'b0100000000;
assign label_9[890] = 10'b0000010000;
assign label_9[891] = 10'b0000000001;
assign label_9[892] = 10'b0100000000;
assign label_9[893] = 10'b0100000000;
assign label_9[894] = 10'b0100000000;
assign label_9[895] = 10'b0100000000;
assign label_9[896] = 10'b0000100000;
assign label_9[897] = 10'b0000100000;
assign label_9[898] = 10'b0000000010;
assign label_9[899] = 10'b0000000010;
assign label_9[900] = 10'b0100000000;
assign label_9[901] = 10'b0100000000;
assign label_9[902] = 10'b0100000000;
assign label_9[903] = 10'b0100000000;
assign label_9[904] = 10'b0100000000;
assign label_9[905] = 10'b0001000000;
assign label_9[906] = 10'b0000000010;
assign label_9[907] = 10'b0001000000;
assign label_9[908] = 10'b0000000100;
assign label_9[909] = 10'b0000000100;
assign label_9[910] = 10'b0001000000;
assign label_9[911] = 10'b0000000100;
assign label_9[912] = 10'b0000000100;
assign label_9[913] = 10'b0001000000;
assign label_9[914] = 10'b0001000000;
assign label_9[915] = 10'b0000000100;
assign label_9[916] = 10'b0000000100;
assign label_9[917] = 10'b0000100000;
assign label_9[918] = 10'b0000000100;
assign label_9[919] = 10'b0000000100;
assign label_9[920] = 10'b0000000010;
assign label_9[921] = 10'b0000100000;
assign label_9[922] = 10'b0000001000;
assign label_9[923] = 10'b0000100000;
assign label_9[924] = 10'b0001000000;
assign label_9[925] = 10'b0001000000;
assign label_9[926] = 10'b0000001000;
assign label_9[927] = 10'b0000001000;
assign label_9[928] = 10'b0001000000;
assign label_9[929] = 10'b0001000000;
assign label_9[930] = 10'b0001000000;
assign label_9[931] = 10'b0000000100;
assign label_9[932] = 10'b0000000100;
assign label_9[933] = 10'b0000000100;
assign label_9[934] = 10'b0000000100;
assign label_9[935] = 10'b0001000000;
assign label_9[936] = 10'b0100000000;
assign label_9[937] = 10'b0001000000;
assign label_9[938] = 10'b0001000000;
assign label_9[939] = 10'b0000100000;
assign label_9[940] = 10'b0100000000;
assign label_9[941] = 10'b0100000000;
assign label_9[942] = 10'b0100000000;
assign label_9[943] = 10'b0000100000;
assign label_9[944] = 10'b0000000100;
assign label_9[945] = 10'b0001000000;
assign label_9[946] = 10'b0000000100;
assign label_9[947] = 10'b0100000000;
assign label_9[948] = 10'b0000000100;
assign label_9[949] = 10'b0100000000;
assign label_9[950] = 10'b0001000000;
assign label_9[951] = 10'b0100000000;
assign label_9[952] = 10'b0000000100;
assign label_9[953] = 10'b0001000000;
assign label_9[954] = 10'b0100000000;
assign label_9[955] = 10'b0000010000;
assign label_9[956] = 10'b0000000100;
assign label_9[957] = 10'b0000000100;
assign label_9[958] = 10'b0100000000;
assign label_9[959] = 10'b1000000000;
assign label_9[960] = 10'b0000000100;
assign label_9[961] = 10'b0000000100;
assign label_9[962] = 10'b0000000100;
assign label_9[963] = 10'b0100000000;
assign label_9[964] = 10'b0001000000;
assign label_9[965] = 10'b0001000000;
assign label_9[966] = 10'b0000000100;
assign label_9[967] = 10'b0000010000;
assign label_9[968] = 10'b0100000000;
assign label_9[969] = 10'b0000000100;
assign label_9[970] = 10'b0000000100;
assign label_9[971] = 10'b0001000000;
assign label_9[972] = 10'b0000000100;
assign label_9[973] = 10'b0100000000;
assign label_9[974] = 10'b0100000000;
assign label_9[975] = 10'b0000000100;
assign label_9[976] = 10'b0100000000;
assign label_9[977] = 10'b0000000010;
assign label_9[978] = 10'b0000000100;
assign label_9[979] = 10'b0000000001;
assign label_9[980] = 10'b0100000000;
assign label_9[981] = 10'b0000000100;
assign label_9[982] = 10'b0001000000;
assign label_9[983] = 10'b0000000001;
assign label_9[984] = 10'b0000010000;
assign label_9[985] = 10'b0000000100;
assign label_9[986] = 10'b0000000100;
assign label_9[987] = 10'b0000000100;
assign label_9[988] = 10'b0000000100;
assign label_9[989] = 10'b0100000000;
assign label_9[990] = 10'b0000000100;
assign label_9[991] = 10'b0000000001;
assign label_9[992] = 10'b0000000100;
assign label_9[993] = 10'b0000000100;
assign label_9[994] = 10'b0000001000;
assign label_9[995] = 10'b0000001000;
assign label_9[996] = 10'b0000000100;
assign label_9[997] = 10'b0000000100;
assign label_9[998] = 10'b0000000010;
assign label_9[999] = 10'b0000000100;
assign label_9[1000] = 10'b0000000100;
assign label_9[1001] = 10'b0000000100;
assign label_9[1002] = 10'b0000000100;
assign label_9[1003] = 10'b0000001000;
assign label_9[1004] = 10'b0000000100;
assign label_9[1005] = 10'b0000000100;
assign label_9[1006] = 10'b0100000000;
assign label_9[1007] = 10'b0000001000;
assign label_9[1008] = 10'b0000000100;
assign label_9[1009] = 10'b0000000100;
assign label_9[1010] = 10'b0000000100;
assign label_9[1011] = 10'b0000000100;
assign label_9[1012] = 10'b0100000000;
assign label_9[1013] = 10'b0000000100;
assign label_9[1014] = 10'b0000000100;
assign label_9[1015] = 10'b0000000100;
assign label_9[1016] = 10'b0000000100;
assign label_9[1017] = 10'b0000000100;
assign label_9[1018] = 10'b0000000100;
assign label_9[1019] = 10'b0000000100;
assign label_9[1020] = 10'b0000001000;
assign label_9[1021] = 10'b0100000000;
assign label_9[1022] = 10'b0000000100;
assign label_9[1023] = 10'b0000000001;
assign feature_index_0[0] = 10'd541;
assign feature_index_0[1] = 10'd403;
assign feature_index_0[2] = 10'd408;
assign feature_index_0[3] = 10'd235;
assign feature_index_0[4] = 10'd652;
assign feature_index_0[5] = 10'd428;
assign feature_index_0[6] = 10'd270;
assign feature_index_0[7] = 10'd457;
assign feature_index_0[8] = 10'd155;
assign feature_index_0[9] = 10'd239;
assign feature_index_0[10] = 10'd319;
assign feature_index_0[11] = 10'd487;
assign feature_index_0[12] = 10'd462;
assign feature_index_0[13] = 10'd683;
assign feature_index_0[14] = 10'd127;
assign feature_index_0[15] = 10'd354;
assign feature_index_0[16] = 10'd97;
assign feature_index_0[17] = 10'd488;
assign feature_index_0[18] = 10'd328;
assign feature_index_0[19] = 10'd71;
assign feature_index_0[20] = 10'd263;
assign feature_index_0[21] = 10'd315;
assign feature_index_0[22] = 10'd328;
assign feature_index_0[23] = 10'd454;
assign feature_index_0[24] = 10'd575;
assign feature_index_0[25] = 10'd626;
assign feature_index_0[26] = 10'd156;
assign feature_index_0[27] = 10'd429;
assign feature_index_0[28] = 10'd466;
assign feature_index_0[29] = 10'd496;
assign feature_index_0[30] = 10'd321;
assign feature_index_0[31] = 10'd461;
assign feature_index_0[32] = 10'd157;
assign feature_index_0[33] = 10'd622;
assign feature_index_0[34] = 10'd511;
assign feature_index_0[35] = 10'd595;
assign feature_index_0[36] = 10'd373;
assign feature_index_0[37] = 10'd455;
assign feature_index_0[38] = 10'd490;
assign feature_index_0[39] = 10'd182;
assign feature_index_0[40] = 10'd0;
assign feature_index_0[41] = 10'd177;
assign feature_index_0[42] = 10'd542;
assign feature_index_0[43] = 10'd483;
assign feature_index_0[44] = 10'd510;
assign feature_index_0[45] = 10'd189;
assign feature_index_0[46] = 10'd510;
assign feature_index_0[47] = 10'd349;
assign feature_index_0[48] = 10'd386;
assign feature_index_0[49] = 10'd653;
assign feature_index_0[50] = 10'd551;
assign feature_index_0[51] = 10'd272;
assign feature_index_0[52] = 10'd290;
assign feature_index_0[53] = 10'd246;
assign feature_index_0[54] = 10'd319;
assign feature_index_0[55] = 10'd490;
assign feature_index_0[56] = 10'd245;
assign feature_index_0[57] = 10'd441;
assign feature_index_0[58] = 10'd513;
assign feature_index_0[59] = 10'd181;
assign feature_index_0[60] = 10'd182;
assign feature_index_0[61] = 10'd488;
assign feature_index_0[62] = 10'd491;
assign feature_index_0[63] = 10'd409;
assign feature_index_0[64] = 10'd495;
assign feature_index_0[65] = 10'd377;
assign feature_index_0[66] = 10'd536;
assign feature_index_0[67] = 10'd265;
assign feature_index_0[68] = 10'd455;
assign feature_index_0[69] = 10'd597;
assign feature_index_0[70] = 10'd425;
assign feature_index_0[71] = 10'd378;
assign feature_index_0[72] = 10'd378;
assign feature_index_0[73] = 10'd398;
assign feature_index_0[74] = 10'd455;
assign feature_index_0[75] = 10'd319;
assign feature_index_0[76] = 10'd461;
assign feature_index_0[77] = 10'd538;
assign feature_index_0[78] = 10'd349;
assign feature_index_0[79] = 10'd97;
assign feature_index_0[80] = 10'd571;
assign feature_index_0[81] = 10'd0;
assign feature_index_0[82] = 10'd0;
assign feature_index_0[83] = 10'd542;
assign feature_index_0[84] = 10'd317;
assign feature_index_0[85] = 10'd298;
assign feature_index_0[86] = 10'd657;
assign feature_index_0[87] = 10'd220;
assign feature_index_0[88] = 10'd374;
assign feature_index_0[89] = 10'd300;
assign feature_index_0[90] = 10'd566;
assign feature_index_0[91] = 10'd578;
assign feature_index_0[92] = 10'd326;
assign feature_index_0[93] = 10'd631;
assign feature_index_0[94] = 10'd412;
assign feature_index_0[95] = 10'd432;
assign feature_index_0[96] = 10'd154;
assign feature_index_0[97] = 10'd342;
assign feature_index_0[98] = 10'd342;
assign feature_index_0[99] = 10'd526;
assign feature_index_0[100] = 10'd182;
assign feature_index_0[101] = 10'd406;
assign feature_index_0[102] = 10'd429;
assign feature_index_0[103] = 10'd241;
assign feature_index_0[104] = 10'd597;
assign feature_index_0[105] = 10'd97;
assign feature_index_0[106] = 10'd379;
assign feature_index_0[107] = 10'd601;
assign feature_index_0[108] = 10'd383;
assign feature_index_0[109] = 10'd661;
assign feature_index_0[110] = 10'd273;
assign feature_index_0[111] = 10'd568;
assign feature_index_0[112] = 10'd296;
assign feature_index_0[113] = 10'd633;
assign feature_index_0[114] = 10'd508;
assign feature_index_0[115] = 10'd665;
assign feature_index_0[116] = 10'd576;
assign feature_index_0[117] = 10'd583;
assign feature_index_0[118] = 10'd355;
assign feature_index_0[119] = 10'd274;
assign feature_index_0[120] = 10'd347;
assign feature_index_0[121] = 10'd386;
assign feature_index_0[122] = 10'd457;
assign feature_index_0[123] = 10'd402;
assign feature_index_0[124] = 10'd318;
assign feature_index_0[125] = 10'd539;
assign feature_index_0[126] = 10'd657;
assign feature_index_0[127] = 10'd399;
assign feature_index_0[128] = 10'd349;
assign feature_index_0[129] = 10'd606;
assign feature_index_0[130] = 10'd633;
assign feature_index_0[131] = 10'd596;
assign feature_index_0[132] = 10'd328;
assign feature_index_0[133] = 10'd516;
assign feature_index_0[134] = 10'd400;
assign feature_index_0[135] = 10'd470;
assign feature_index_0[136] = 10'd286;
assign feature_index_0[137] = 10'd186;
assign feature_index_0[138] = 10'd652;
assign feature_index_0[139] = 10'd470;
assign feature_index_0[140] = 10'd0;
assign feature_index_0[141] = 10'd0;
assign feature_index_0[142] = 10'd0;
assign feature_index_0[143] = 10'd459;
assign feature_index_0[144] = 10'd183;
assign feature_index_0[145] = 10'd353;
assign feature_index_0[146] = 10'd299;
assign feature_index_0[147] = 10'd582;
assign feature_index_0[148] = 10'd191;
assign feature_index_0[149] = 10'd69;
assign feature_index_0[150] = 10'd237;
assign feature_index_0[151] = 10'd489;
assign feature_index_0[152] = 10'd297;
assign feature_index_0[153] = 10'd653;
assign feature_index_0[154] = 10'd574;
assign feature_index_0[155] = 10'd622;
assign feature_index_0[156] = 10'd408;
assign feature_index_0[157] = 10'd372;
assign feature_index_0[158] = 10'd694;
assign feature_index_0[159] = 10'd526;
assign feature_index_0[160] = 10'd597;
assign feature_index_0[161] = 10'd626;
assign feature_index_0[162] = 10'd100;
assign feature_index_0[163] = 10'd0;
assign feature_index_0[164] = 10'd0;
assign feature_index_0[165] = 10'd0;
assign feature_index_0[166] = 10'd0;
assign feature_index_0[167] = 10'd568;
assign feature_index_0[168] = 10'd242;
assign feature_index_0[169] = 10'd659;
assign feature_index_0[170] = 10'd599;
assign feature_index_0[171] = 10'd355;
assign feature_index_0[172] = 10'd151;
assign feature_index_0[173] = 10'd375;
assign feature_index_0[174] = 10'd550;
assign feature_index_0[175] = 10'd182;
assign feature_index_0[176] = 10'd209;
assign feature_index_0[177] = 10'd129;
assign feature_index_0[178] = 10'd351;
assign feature_index_0[179] = 10'd540;
assign feature_index_0[180] = 10'd185;
assign feature_index_0[181] = 10'd0;
assign feature_index_0[182] = 10'd292;
assign feature_index_0[183] = 10'd181;
assign feature_index_0[184] = 10'd325;
assign feature_index_0[185] = 10'd331;
assign feature_index_0[186] = 10'd272;
assign feature_index_0[187] = 10'd709;
assign feature_index_0[188] = 10'd324;
assign feature_index_0[189] = 10'd379;
assign feature_index_0[190] = 10'd433;
assign feature_index_0[191] = 10'd566;
assign feature_index_0[192] = 10'd413;
assign feature_index_0[193] = 10'd539;
assign feature_index_0[194] = 10'd462;
assign feature_index_0[195] = 10'd154;
assign feature_index_0[196] = 10'd519;
assign feature_index_0[197] = 10'd343;
assign feature_index_0[198] = 10'd461;
assign feature_index_0[199] = 10'd180;
assign feature_index_0[200] = 10'd609;
assign feature_index_0[201] = 10'd579;
assign feature_index_0[202] = 10'd380;
assign feature_index_0[203] = 10'd656;
assign feature_index_0[204] = 10'd607;
assign feature_index_0[205] = 10'd359;
assign feature_index_0[206] = 10'd483;
assign feature_index_0[207] = 10'd173;
assign feature_index_0[208] = 10'd582;
assign feature_index_0[209] = 10'd326;
assign feature_index_0[210] = 10'd407;
assign feature_index_0[211] = 10'd272;
assign feature_index_0[212] = 10'd517;
assign feature_index_0[213] = 10'd357;
assign feature_index_0[214] = 10'd268;
assign feature_index_0[215] = 10'd606;
assign feature_index_0[216] = 10'd183;
assign feature_index_0[217] = 10'd360;
assign feature_index_0[218] = 10'd266;
assign feature_index_0[219] = 10'd509;
assign feature_index_0[220] = 10'd328;
assign feature_index_0[221] = 10'd243;
assign feature_index_0[222] = 10'd385;
assign feature_index_0[223] = 10'd655;
assign feature_index_0[224] = 10'd326;
assign feature_index_0[225] = 10'd399;
assign feature_index_0[226] = 10'd186;
assign feature_index_0[227] = 10'd602;
assign feature_index_0[228] = 10'd657;
assign feature_index_0[229] = 10'd300;
assign feature_index_0[230] = 10'd372;
assign feature_index_0[231] = 10'd691;
assign feature_index_0[232] = 10'd0;
assign feature_index_0[233] = 10'd527;
assign feature_index_0[234] = 10'd485;
assign feature_index_0[235] = 10'd355;
assign feature_index_0[236] = 10'd0;
assign feature_index_0[237] = 10'd299;
assign feature_index_0[238] = 10'd186;
assign feature_index_0[239] = 10'd575;
assign feature_index_0[240] = 10'd212;
assign feature_index_0[241] = 10'd580;
assign feature_index_0[242] = 10'd376;
assign feature_index_0[243] = 10'd489;
assign feature_index_0[244] = 10'd570;
assign feature_index_0[245] = 10'd520;
assign feature_index_0[246] = 10'd660;
assign feature_index_0[247] = 10'd630;
assign feature_index_0[248] = 10'd518;
assign feature_index_0[249] = 10'd316;
assign feature_index_0[250] = 10'd540;
assign feature_index_0[251] = 10'd514;
assign feature_index_0[252] = 10'd430;
assign feature_index_0[253] = 10'd525;
assign feature_index_0[254] = 10'd410;
assign feature_index_0[255] = 10'd328;
assign feature_index_0[256] = 10'd598;
assign feature_index_0[257] = 10'd318;
assign feature_index_0[258] = 10'd288;
assign feature_index_0[259] = 10'd316;
assign feature_index_0[260] = 10'd236;
assign feature_index_0[261] = 10'd527;
assign feature_index_0[262] = 10'd346;
assign feature_index_0[263] = 10'd211;
assign feature_index_0[264] = 10'd708;
assign feature_index_0[265] = 10'd182;
assign feature_index_0[266] = 10'd185;
assign feature_index_0[267] = 10'd134;
assign feature_index_0[268] = 10'd178;
assign feature_index_0[269] = 10'd213;
assign feature_index_0[270] = 10'd324;
assign feature_index_0[271] = 10'd568;
assign feature_index_0[272] = 10'd526;
assign feature_index_0[273] = 10'd382;
assign feature_index_0[274] = 10'd348;
assign feature_index_0[275] = 10'd0;
assign feature_index_0[276] = 10'd296;
assign feature_index_0[277] = 10'd320;
assign feature_index_0[278] = 10'd372;
assign feature_index_0[279] = 10'd261;
assign feature_index_0[280] = 10'd372;
assign feature_index_0[281] = 10'd0;
assign feature_index_0[282] = 10'd0;
assign feature_index_0[283] = 10'd0;
assign feature_index_0[284] = 10'd0;
assign feature_index_0[285] = 10'd0;
assign feature_index_0[286] = 10'd0;
assign feature_index_0[287] = 10'd148;
assign feature_index_0[288] = 10'd483;
assign feature_index_0[289] = 10'd286;
assign feature_index_0[290] = 10'd345;
assign feature_index_0[291] = 10'd437;
assign feature_index_0[292] = 10'd274;
assign feature_index_0[293] = 10'd173;
assign feature_index_0[294] = 10'd290;
assign feature_index_0[295] = 10'd348;
assign feature_index_0[296] = 10'd680;
assign feature_index_0[297] = 10'd210;
assign feature_index_0[298] = 10'd213;
assign feature_index_0[299] = 10'd239;
assign feature_index_0[300] = 10'd0;
assign feature_index_0[301] = 10'd124;
assign feature_index_0[302] = 10'd347;
assign feature_index_0[303] = 10'd219;
assign feature_index_0[304] = 10'd404;
assign feature_index_0[305] = 10'd579;
assign feature_index_0[306] = 10'd411;
assign feature_index_0[307] = 10'd262;
assign feature_index_0[308] = 10'd431;
assign feature_index_0[309] = 10'd442;
assign feature_index_0[310] = 10'd572;
assign feature_index_0[311] = 10'd356;
assign feature_index_0[312] = 10'd406;
assign feature_index_0[313] = 10'd382;
assign feature_index_0[314] = 10'd376;
assign feature_index_0[315] = 10'd573;
assign feature_index_0[316] = 10'd626;
assign feature_index_0[317] = 10'd462;
assign feature_index_0[318] = 10'd0;
assign feature_index_0[319] = 10'd400;
assign feature_index_0[320] = 10'd694;
assign feature_index_0[321] = 10'd425;
assign feature_index_0[322] = 10'd296;
assign feature_index_0[323] = 10'd273;
assign feature_index_0[324] = 10'd491;
assign feature_index_0[325] = 10'd411;
assign feature_index_0[326] = 10'd301;
assign feature_index_0[327] = 10'd0;
assign feature_index_0[328] = 10'd0;
assign feature_index_0[329] = 10'd0;
assign feature_index_0[330] = 10'd0;
assign feature_index_0[331] = 10'd0;
assign feature_index_0[332] = 10'd0;
assign feature_index_0[333] = 10'd0;
assign feature_index_0[334] = 10'd0;
assign feature_index_0[335] = 10'd181;
assign feature_index_0[336] = 10'd381;
assign feature_index_0[337] = 10'd466;
assign feature_index_0[338] = 10'd545;
assign feature_index_0[339] = 10'd260;
assign feature_index_0[340] = 10'd372;
assign feature_index_0[341] = 10'd344;
assign feature_index_0[342] = 10'd272;
assign feature_index_0[343] = 10'd627;
assign feature_index_0[344] = 10'd348;
assign feature_index_0[345] = 10'd539;
assign feature_index_0[346] = 10'd181;
assign feature_index_0[347] = 10'd298;
assign feature_index_0[348] = 10'd299;
assign feature_index_0[349] = 10'd656;
assign feature_index_0[350] = 10'd460;
assign feature_index_0[351] = 10'd191;
assign feature_index_0[352] = 10'd325;
assign feature_index_0[353] = 10'd0;
assign feature_index_0[354] = 10'd599;
assign feature_index_0[355] = 10'd350;
assign feature_index_0[356] = 10'd296;
assign feature_index_0[357] = 10'd218;
assign feature_index_0[358] = 10'd545;
assign feature_index_0[359] = 10'd191;
assign feature_index_0[360] = 10'd351;
assign feature_index_0[361] = 10'd270;
assign feature_index_0[362] = 10'd542;
assign feature_index_0[363] = 10'd0;
assign feature_index_0[364] = 10'd0;
assign feature_index_0[365] = 10'd185;
assign feature_index_0[366] = 10'd296;
assign feature_index_0[367] = 10'd481;
assign feature_index_0[368] = 10'd262;
assign feature_index_0[369] = 10'd296;
assign feature_index_0[370] = 10'd274;
assign feature_index_0[371] = 10'd264;
assign feature_index_0[372] = 10'd355;
assign feature_index_0[373] = 10'd630;
assign feature_index_0[374] = 10'd516;
assign feature_index_0[375] = 10'd192;
assign feature_index_0[376] = 10'd187;
assign feature_index_0[377] = 10'd571;
assign feature_index_0[378] = 10'd289;
assign feature_index_0[379] = 10'd276;
assign feature_index_0[380] = 10'd457;
assign feature_index_0[381] = 10'd205;
assign feature_index_0[382] = 10'd519;
assign feature_index_0[383] = 10'd485;
assign feature_index_0[384] = 10'd398;
assign feature_index_0[385] = 10'd149;
assign feature_index_0[386] = 10'd347;
assign feature_index_0[387] = 10'd326;
assign feature_index_0[388] = 10'd176;
assign feature_index_0[389] = 10'd290;
assign feature_index_0[390] = 10'd71;
assign feature_index_0[391] = 10'd321;
assign feature_index_0[392] = 10'd290;
assign feature_index_0[393] = 10'd417;
assign feature_index_0[394] = 10'd359;
assign feature_index_0[395] = 10'd152;
assign feature_index_0[396] = 10'd0;
assign feature_index_0[397] = 10'd70;
assign feature_index_0[398] = 10'd0;
assign feature_index_0[399] = 10'd324;
assign feature_index_0[400] = 10'd540;
assign feature_index_0[401] = 10'd521;
assign feature_index_0[402] = 10'd579;
assign feature_index_0[403] = 10'd512;
assign feature_index_0[404] = 10'd377;
assign feature_index_0[405] = 10'd651;
assign feature_index_0[406] = 10'd466;
assign feature_index_0[407] = 10'd403;
assign feature_index_0[408] = 10'd376;
assign feature_index_0[409] = 10'd438;
assign feature_index_0[410] = 10'd660;
assign feature_index_0[411] = 10'd347;
assign feature_index_0[412] = 10'd377;
assign feature_index_0[413] = 10'd554;
assign feature_index_0[414] = 10'd552;
assign feature_index_0[415] = 10'd369;
assign feature_index_0[416] = 10'd0;
assign feature_index_0[417] = 10'd378;
assign feature_index_0[418] = 10'd375;
assign feature_index_0[419] = 10'd598;
assign feature_index_0[420] = 10'd216;
assign feature_index_0[421] = 10'd292;
assign feature_index_0[422] = 10'd274;
assign feature_index_0[423] = 10'd484;
assign feature_index_0[424] = 10'd379;
assign feature_index_0[425] = 10'd103;
assign feature_index_0[426] = 10'd188;
assign feature_index_0[427] = 10'd221;
assign feature_index_0[428] = 10'd352;
assign feature_index_0[429] = 10'd242;
assign feature_index_0[430] = 10'd146;
assign feature_index_0[431] = 10'd400;
assign feature_index_0[432] = 10'd437;
assign feature_index_0[433] = 10'd218;
assign feature_index_0[434] = 10'd125;
assign feature_index_0[435] = 10'd352;
assign feature_index_0[436] = 10'd686;
assign feature_index_0[437] = 10'd376;
assign feature_index_0[438] = 10'd711;
assign feature_index_0[439] = 10'd431;
assign feature_index_0[440] = 10'd0;
assign feature_index_0[441] = 10'd352;
assign feature_index_0[442] = 10'd398;
assign feature_index_0[443] = 10'd289;
assign feature_index_0[444] = 10'd94;
assign feature_index_0[445] = 10'd134;
assign feature_index_0[446] = 10'd602;
assign feature_index_0[447] = 10'd206;
assign feature_index_0[448] = 10'd405;
assign feature_index_0[449] = 10'd386;
assign feature_index_0[450] = 10'd437;
assign feature_index_0[451] = 10'd658;
assign feature_index_0[452] = 10'd188;
assign feature_index_0[453] = 10'd400;
assign feature_index_0[454] = 10'd189;
assign feature_index_0[455] = 10'd501;
assign feature_index_0[456] = 10'd637;
assign feature_index_0[457] = 10'd630;
assign feature_index_0[458] = 10'd176;
assign feature_index_0[459] = 10'd156;
assign feature_index_0[460] = 10'd157;
assign feature_index_0[461] = 10'd552;
assign feature_index_0[462] = 10'd343;
assign feature_index_0[463] = 10'd635;
assign feature_index_0[464] = 10'd0;
assign feature_index_0[465] = 10'd0;
assign feature_index_0[466] = 10'd0;
assign feature_index_0[467] = 10'd0;
assign feature_index_0[468] = 10'd0;
assign feature_index_0[469] = 10'd0;
assign feature_index_0[470] = 10'd433;
assign feature_index_0[471] = 10'd158;
assign feature_index_0[472] = 10'd435;
assign feature_index_0[473] = 10'd0;
assign feature_index_0[474] = 10'd0;
assign feature_index_0[475] = 10'd488;
assign feature_index_0[476] = 10'd0;
assign feature_index_0[477] = 10'd0;
assign feature_index_0[478] = 10'd156;
assign feature_index_0[479] = 10'd373;
assign feature_index_0[480] = 10'd439;
assign feature_index_0[481] = 10'd187;
assign feature_index_0[482] = 10'd432;
assign feature_index_0[483] = 10'd316;
assign feature_index_0[484] = 10'd373;
assign feature_index_0[485] = 10'd485;
assign feature_index_0[486] = 10'd462;
assign feature_index_0[487] = 10'd598;
assign feature_index_0[488] = 10'd344;
assign feature_index_0[489] = 10'd637;
assign feature_index_0[490] = 10'd238;
assign feature_index_0[491] = 10'd296;
assign feature_index_0[492] = 10'd684;
assign feature_index_0[493] = 10'd526;
assign feature_index_0[494] = 10'd657;
assign feature_index_0[495] = 10'd159;
assign feature_index_0[496] = 10'd406;
assign feature_index_0[497] = 10'd406;
assign feature_index_0[498] = 10'd318;
assign feature_index_0[499] = 10'd656;
assign feature_index_0[500] = 10'd575;
assign feature_index_0[501] = 10'd431;
assign feature_index_0[502] = 10'd659;
assign feature_index_0[503] = 10'd484;
assign feature_index_0[504] = 10'd269;
assign feature_index_0[505] = 10'd296;
assign feature_index_0[506] = 10'd374;
assign feature_index_0[507] = 10'd235;
assign feature_index_0[508] = 10'd351;
assign feature_index_0[509] = 10'd319;
assign feature_index_0[510] = 10'd399;
assign feature_index_0[511] = 10'd522;
assign feature_index_0[512] = 10'd567;
assign feature_index_0[513] = 10'd566;
assign feature_index_0[514] = 10'd535;
assign feature_index_0[515] = 10'd404;
assign feature_index_0[516] = 10'd125;
assign feature_index_0[517] = 10'd265;
assign feature_index_0[518] = 10'd268;
assign feature_index_0[519] = 10'd438;
assign feature_index_0[520] = 10'd210;
assign feature_index_0[521] = 10'd318;
assign feature_index_0[522] = 10'd491;
assign feature_index_0[523] = 10'd215;
assign feature_index_0[524] = 10'd0;
assign feature_index_0[525] = 10'd261;
assign feature_index_0[526] = 10'd624;
assign feature_index_0[527] = 10'd513;
assign feature_index_0[528] = 10'd155;
assign feature_index_0[529] = 10'd183;
assign feature_index_0[530] = 10'd0;
assign feature_index_0[531] = 10'd604;
assign feature_index_0[532] = 10'd655;
assign feature_index_0[533] = 10'd406;
assign feature_index_0[534] = 10'd465;
assign feature_index_0[535] = 10'd554;
assign feature_index_0[536] = 10'd302;
assign feature_index_0[537] = 10'd297;
assign feature_index_0[538] = 10'd432;
assign feature_index_0[539] = 10'd517;
assign feature_index_0[540] = 10'd0;
assign feature_index_0[541] = 10'd0;
assign feature_index_0[542] = 10'd567;
assign feature_index_0[543] = 10'd437;
assign feature_index_0[544] = 10'd320;
assign feature_index_0[545] = 10'd486;
assign feature_index_0[546] = 10'd577;
assign feature_index_0[547] = 10'd595;
assign feature_index_0[548] = 10'd739;
assign feature_index_0[549] = 10'd452;
assign feature_index_0[550] = 10'd0;
assign feature_index_0[551] = 10'd0;
assign feature_index_0[552] = 10'd0;
assign feature_index_0[553] = 10'd680;
assign feature_index_0[554] = 10'd193;
assign feature_index_0[555] = 10'd0;
assign feature_index_0[556] = 10'd236;
assign feature_index_0[557] = 10'd128;
assign feature_index_0[558] = 10'd404;
assign feature_index_0[559] = 10'd0;
assign feature_index_0[560] = 10'd155;
assign feature_index_0[561] = 10'd0;
assign feature_index_0[562] = 10'd0;
assign feature_index_0[563] = 10'd0;
assign feature_index_0[564] = 10'd0;
assign feature_index_0[565] = 10'd0;
assign feature_index_0[566] = 10'd0;
assign feature_index_0[567] = 10'd0;
assign feature_index_0[568] = 10'd0;
assign feature_index_0[569] = 10'd0;
assign feature_index_0[570] = 10'd0;
assign feature_index_0[571] = 10'd0;
assign feature_index_0[572] = 10'd0;
assign feature_index_0[573] = 10'd0;
assign feature_index_0[574] = 10'd0;
assign feature_index_0[575] = 10'd514;
assign feature_index_0[576] = 10'd210;
assign feature_index_0[577] = 10'd160;
assign feature_index_0[578] = 10'd184;
assign feature_index_0[579] = 10'd232;
assign feature_index_0[580] = 10'd515;
assign feature_index_0[581] = 10'd376;
assign feature_index_0[582] = 10'd326;
assign feature_index_0[583] = 10'd146;
assign feature_index_0[584] = 10'd706;
assign feature_index_0[585] = 10'd208;
assign feature_index_0[586] = 10'd216;
assign feature_index_0[587] = 10'd470;
assign feature_index_0[588] = 10'd0;
assign feature_index_0[589] = 10'd206;
assign feature_index_0[590] = 10'd528;
assign feature_index_0[591] = 10'd344;
assign feature_index_0[592] = 10'd153;
assign feature_index_0[593] = 10'd572;
assign feature_index_0[594] = 10'd0;
assign feature_index_0[595] = 10'd231;
assign feature_index_0[596] = 10'd370;
assign feature_index_0[597] = 10'd0;
assign feature_index_0[598] = 10'd573;
assign feature_index_0[599] = 10'd210;
assign feature_index_0[600] = 10'd457;
assign feature_index_0[601] = 10'd0;
assign feature_index_0[602] = 10'd0;
assign feature_index_0[603] = 10'd717;
assign feature_index_0[604] = 10'd300;
assign feature_index_0[605] = 10'd238;
assign feature_index_0[606] = 10'd267;
assign feature_index_0[607] = 10'd351;
assign feature_index_0[608] = 10'd662;
assign feature_index_0[609] = 10'd349;
assign feature_index_0[610] = 10'd298;
assign feature_index_0[611] = 10'd323;
assign feature_index_0[612] = 10'd268;
assign feature_index_0[613] = 10'd649;
assign feature_index_0[614] = 10'd460;
assign feature_index_0[615] = 10'd0;
assign feature_index_0[616] = 10'd288;
assign feature_index_0[617] = 10'd303;
assign feature_index_0[618] = 10'd0;
assign feature_index_0[619] = 10'd382;
assign feature_index_0[620] = 10'd412;
assign feature_index_0[621] = 10'd435;
assign feature_index_0[622] = 10'd294;
assign feature_index_0[623] = 10'd412;
assign feature_index_0[624] = 10'd159;
assign feature_index_0[625] = 10'd291;
assign feature_index_0[626] = 10'd0;
assign feature_index_0[627] = 10'd201;
assign feature_index_0[628] = 10'd376;
assign feature_index_0[629] = 10'd370;
assign feature_index_0[630] = 10'd330;
assign feature_index_0[631] = 10'd460;
assign feature_index_0[632] = 10'd654;
assign feature_index_0[633] = 10'd486;
assign feature_index_0[634] = 10'd567;
assign feature_index_0[635] = 10'd0;
assign feature_index_0[636] = 10'd158;
assign feature_index_0[637] = 10'd0;
assign feature_index_0[638] = 10'd0;
assign feature_index_0[639] = 10'd436;
assign feature_index_0[640] = 10'd294;
assign feature_index_0[641] = 10'd455;
assign feature_index_0[642] = 10'd294;
assign feature_index_0[643] = 10'd509;
assign feature_index_0[644] = 10'd0;
assign feature_index_0[645] = 10'd430;
assign feature_index_0[646] = 10'd211;
assign feature_index_0[647] = 10'd212;
assign feature_index_0[648] = 10'd212;
assign feature_index_0[649] = 10'd345;
assign feature_index_0[650] = 10'd150;
assign feature_index_0[651] = 10'd298;
assign feature_index_0[652] = 10'd544;
assign feature_index_0[653] = 10'd325;
assign feature_index_0[654] = 10'd0;
assign feature_index_0[655] = 10'd0;
assign feature_index_0[656] = 10'd0;
assign feature_index_0[657] = 10'd0;
assign feature_index_0[658] = 10'd0;
assign feature_index_0[659] = 10'd0;
assign feature_index_0[660] = 10'd0;
assign feature_index_0[661] = 10'd0;
assign feature_index_0[662] = 10'd0;
assign feature_index_0[663] = 10'd0;
assign feature_index_0[664] = 10'd0;
assign feature_index_0[665] = 10'd0;
assign feature_index_0[666] = 10'd0;
assign feature_index_0[667] = 10'd0;
assign feature_index_0[668] = 10'd0;
assign feature_index_0[669] = 10'd0;
assign feature_index_0[670] = 10'd0;
assign feature_index_0[671] = 10'd101;
assign feature_index_0[672] = 10'd373;
assign feature_index_0[673] = 10'd462;
assign feature_index_0[674] = 10'd577;
assign feature_index_0[675] = 10'd157;
assign feature_index_0[676] = 10'd96;
assign feature_index_0[677] = 10'd124;
assign feature_index_0[678] = 10'd594;
assign feature_index_0[679] = 10'd485;
assign feature_index_0[680] = 10'd516;
assign feature_index_0[681] = 10'd119;
assign feature_index_0[682] = 10'd314;
assign feature_index_0[683] = 10'd373;
assign feature_index_0[684] = 10'd235;
assign feature_index_0[685] = 10'd468;
assign feature_index_0[686] = 10'd259;
assign feature_index_0[687] = 10'd352;
assign feature_index_0[688] = 10'd323;
assign feature_index_0[689] = 10'd564;
assign feature_index_0[690] = 10'd465;
assign feature_index_0[691] = 10'd516;
assign feature_index_0[692] = 10'd374;
assign feature_index_0[693] = 10'd609;
assign feature_index_0[694] = 10'd317;
assign feature_index_0[695] = 10'd414;
assign feature_index_0[696] = 10'd343;
assign feature_index_0[697] = 10'd549;
assign feature_index_0[698] = 10'd718;
assign feature_index_0[699] = 10'd573;
assign feature_index_0[700] = 10'd414;
assign feature_index_0[701] = 10'd289;
assign feature_index_0[702] = 10'd293;
assign feature_index_0[703] = 10'd680;
assign feature_index_0[704] = 10'd134;
assign feature_index_0[705] = 10'd269;
assign feature_index_0[706] = 10'd518;
assign feature_index_0[707] = 10'd0;
assign feature_index_0[708] = 10'd0;
assign feature_index_0[709] = 10'd0;
assign feature_index_0[710] = 10'd679;
assign feature_index_0[711] = 10'd150;
assign feature_index_0[712] = 10'd164;
assign feature_index_0[713] = 10'd462;
assign feature_index_0[714] = 10'd456;
assign feature_index_0[715] = 10'd681;
assign feature_index_0[716] = 10'd244;
assign feature_index_0[717] = 10'd134;
assign feature_index_0[718] = 10'd548;
assign feature_index_0[719] = 10'd353;
assign feature_index_0[720] = 10'd0;
assign feature_index_0[721] = 10'd0;
assign feature_index_0[722] = 10'd233;
assign feature_index_0[723] = 10'd0;
assign feature_index_0[724] = 10'd353;
assign feature_index_0[725] = 10'd511;
assign feature_index_0[726] = 10'd678;
assign feature_index_0[727] = 10'd0;
assign feature_index_0[728] = 10'd0;
assign feature_index_0[729] = 10'd0;
assign feature_index_0[730] = 10'd0;
assign feature_index_0[731] = 10'd0;
assign feature_index_0[732] = 10'd528;
assign feature_index_0[733] = 10'd0;
assign feature_index_0[734] = 10'd0;
assign feature_index_0[735] = 10'd325;
assign feature_index_0[736] = 10'd409;
assign feature_index_0[737] = 10'd206;
assign feature_index_0[738] = 10'd273;
assign feature_index_0[739] = 10'd236;
assign feature_index_0[740] = 10'd348;
assign feature_index_0[741] = 10'd271;
assign feature_index_0[742] = 10'd330;
assign feature_index_0[743] = 10'd299;
assign feature_index_0[744] = 10'd537;
assign feature_index_0[745] = 10'd437;
assign feature_index_0[746] = 10'd0;
assign feature_index_0[747] = 10'd628;
assign feature_index_0[748] = 10'd351;
assign feature_index_0[749] = 10'd289;
assign feature_index_0[750] = 10'd275;
assign feature_index_0[751] = 10'd381;
assign feature_index_0[752] = 10'd538;
assign feature_index_0[753] = 10'd232;
assign feature_index_0[754] = 10'd675;
assign feature_index_0[755] = 10'd235;
assign feature_index_0[756] = 10'd429;
assign feature_index_0[757] = 10'd523;
assign feature_index_0[758] = 10'd428;
assign feature_index_0[759] = 10'd597;
assign feature_index_0[760] = 10'd650;
assign feature_index_0[761] = 10'd303;
assign feature_index_0[762] = 10'd0;
assign feature_index_0[763] = 10'd548;
assign feature_index_0[764] = 10'd295;
assign feature_index_0[765] = 10'd563;
assign feature_index_0[766] = 10'd490;
assign feature_index_0[767] = 10'd327;
assign feature_index_0[768] = 10'd627;
assign feature_index_0[769] = 10'd657;
assign feature_index_0[770] = 10'd128;
assign feature_index_0[771] = 10'd379;
assign feature_index_0[772] = 10'd0;
assign feature_index_0[773] = 10'd0;
assign feature_index_0[774] = 10'd0;
assign feature_index_0[775] = 10'd246;
assign feature_index_0[776] = 10'd600;
assign feature_index_0[777] = 10'd491;
assign feature_index_0[778] = 10'd467;
assign feature_index_0[779] = 10'd322;
assign feature_index_0[780] = 10'd126;
assign feature_index_0[781] = 10'd265;
assign feature_index_0[782] = 10'd0;
assign feature_index_0[783] = 10'd0;
assign feature_index_0[784] = 10'd424;
assign feature_index_0[785] = 10'd436;
assign feature_index_0[786] = 10'd464;
assign feature_index_0[787] = 10'd0;
assign feature_index_0[788] = 10'd0;
assign feature_index_0[789] = 10'd0;
assign feature_index_0[790] = 10'd0;
assign feature_index_0[791] = 10'd239;
assign feature_index_0[792] = 10'd331;
assign feature_index_0[793] = 10'd0;
assign feature_index_0[794] = 10'd0;
assign feature_index_0[795] = 10'd245;
assign feature_index_0[796] = 10'd0;
assign feature_index_0[797] = 10'd0;
assign feature_index_0[798] = 10'd0;
assign feature_index_0[799] = 10'd357;
assign feature_index_0[800] = 10'd304;
assign feature_index_0[801] = 10'd378;
assign feature_index_0[802] = 10'd688;
assign feature_index_0[803] = 10'd460;
assign feature_index_0[804] = 10'd0;
assign feature_index_0[805] = 10'd491;
assign feature_index_0[806] = 10'd153;
assign feature_index_0[807] = 10'd135;
assign feature_index_0[808] = 10'd403;
assign feature_index_0[809] = 10'd274;
assign feature_index_0[810] = 10'd0;
assign feature_index_0[811] = 10'd464;
assign feature_index_0[812] = 10'd436;
assign feature_index_0[813] = 10'd579;
assign feature_index_0[814] = 10'd273;
assign feature_index_0[815] = 10'd455;
assign feature_index_0[816] = 10'd125;
assign feature_index_0[817] = 10'd125;
assign feature_index_0[818] = 10'd190;
assign feature_index_0[819] = 10'd240;
assign feature_index_0[820] = 10'd299;
assign feature_index_0[821] = 10'd0;
assign feature_index_0[822] = 10'd491;
assign feature_index_0[823] = 10'd190;
assign feature_index_0[824] = 10'd382;
assign feature_index_0[825] = 10'd411;
assign feature_index_0[826] = 10'd302;
assign feature_index_0[827] = 10'd658;
assign feature_index_0[828] = 10'd464;
assign feature_index_0[829] = 10'd245;
assign feature_index_0[830] = 10'd0;
assign feature_index_0[831] = 10'd248;
assign feature_index_0[832] = 10'd202;
assign feature_index_0[833] = 10'd0;
assign feature_index_0[834] = 10'd0;
assign feature_index_0[835] = 10'd102;
assign feature_index_0[836] = 10'd438;
assign feature_index_0[837] = 10'd0;
assign feature_index_0[838] = 10'd382;
assign feature_index_0[839] = 10'd544;
assign feature_index_0[840] = 10'd461;
assign feature_index_0[841] = 10'd210;
assign feature_index_0[842] = 10'd354;
assign feature_index_0[843] = 10'd442;
assign feature_index_0[844] = 10'd648;
assign feature_index_0[845] = 10'd0;
assign feature_index_0[846] = 10'd0;
assign feature_index_0[847] = 10'd127;
assign feature_index_0[848] = 10'd405;
assign feature_index_0[849] = 10'd628;
assign feature_index_0[850] = 10'd414;
assign feature_index_0[851] = 10'd130;
assign feature_index_0[852] = 10'd404;
assign feature_index_0[853] = 10'd0;
assign feature_index_0[854] = 10'd315;
assign feature_index_0[855] = 10'd99;
assign feature_index_0[856] = 10'd0;
assign feature_index_0[857] = 10'd568;
assign feature_index_0[858] = 10'd101;
assign feature_index_0[859] = 10'd327;
assign feature_index_0[860] = 10'd353;
assign feature_index_0[861] = 10'd373;
assign feature_index_0[862] = 10'd239;
assign feature_index_0[863] = 10'd245;
assign feature_index_0[864] = 10'd345;
assign feature_index_0[865] = 10'd465;
assign feature_index_0[866] = 10'd658;
assign feature_index_0[867] = 10'd368;
assign feature_index_0[868] = 10'd159;
assign feature_index_0[869] = 10'd318;
assign feature_index_0[870] = 10'd241;
assign feature_index_0[871] = 10'd331;
assign feature_index_0[872] = 10'd304;
assign feature_index_0[873] = 10'd0;
assign feature_index_0[874] = 10'd0;
assign feature_index_0[875] = 10'd269;
assign feature_index_0[876] = 10'd495;
assign feature_index_0[877] = 10'd400;
assign feature_index_0[878] = 10'd456;
assign feature_index_0[879] = 10'd570;
assign feature_index_0[880] = 10'd662;
assign feature_index_0[881] = 10'd0;
assign feature_index_0[882] = 10'd0;
assign feature_index_0[883] = 10'd374;
assign feature_index_0[884] = 10'd268;
assign feature_index_0[885] = 10'd0;
assign feature_index_0[886] = 10'd245;
assign feature_index_0[887] = 10'd465;
assign feature_index_0[888] = 10'd192;
assign feature_index_0[889] = 10'd316;
assign feature_index_0[890] = 10'd0;
assign feature_index_0[891] = 10'd379;
assign feature_index_0[892] = 10'd0;
assign feature_index_0[893] = 10'd548;
assign feature_index_0[894] = 10'd321;
assign feature_index_0[895] = 10'd245;
assign feature_index_0[896] = 10'd631;
assign feature_index_0[897] = 10'd239;
assign feature_index_0[898] = 10'd326;
assign feature_index_0[899] = 10'd235;
assign feature_index_0[900] = 10'd272;
assign feature_index_0[901] = 10'd206;
assign feature_index_0[902] = 10'd457;
assign feature_index_0[903] = 10'd653;
assign feature_index_0[904] = 10'd369;
assign feature_index_0[905] = 10'd243;
assign feature_index_0[906] = 10'd162;
assign feature_index_0[907] = 10'd149;
assign feature_index_0[908] = 10'd180;
assign feature_index_0[909] = 10'd494;
assign feature_index_0[910] = 10'd653;
assign feature_index_0[911] = 10'd573;
assign feature_index_0[912] = 10'd240;
assign feature_index_0[913] = 10'd162;
assign feature_index_0[914] = 10'd608;
assign feature_index_0[915] = 10'd400;
assign feature_index_0[916] = 10'd269;
assign feature_index_0[917] = 10'd353;
assign feature_index_0[918] = 10'd288;
assign feature_index_0[919] = 10'd273;
assign feature_index_0[920] = 10'd653;
assign feature_index_0[921] = 10'd427;
assign feature_index_0[922] = 10'd655;
assign feature_index_0[923] = 10'd273;
assign feature_index_0[924] = 10'd0;
assign feature_index_0[925] = 10'd451;
assign feature_index_0[926] = 10'd157;
assign feature_index_0[927] = 10'd486;
assign feature_index_0[928] = 10'd401;
assign feature_index_0[929] = 10'd0;
assign feature_index_0[930] = 10'd0;
assign feature_index_0[931] = 10'd0;
assign feature_index_0[932] = 10'd0;
assign feature_index_0[933] = 10'd0;
assign feature_index_0[934] = 10'd0;
assign feature_index_0[935] = 10'd0;
assign feature_index_0[936] = 10'd0;
assign feature_index_0[937] = 10'd0;
assign feature_index_0[938] = 10'd0;
assign feature_index_0[939] = 10'd0;
assign feature_index_0[940] = 10'd0;
assign feature_index_0[941] = 10'd0;
assign feature_index_0[942] = 10'd0;
assign feature_index_0[943] = 10'd433;
assign feature_index_0[944] = 10'd633;
assign feature_index_0[945] = 10'd188;
assign feature_index_0[946] = 10'd0;
assign feature_index_0[947] = 10'd0;
assign feature_index_0[948] = 10'd0;
assign feature_index_0[949] = 10'd0;
assign feature_index_0[950] = 10'd0;
assign feature_index_0[951] = 10'd187;
assign feature_index_0[952] = 10'd374;
assign feature_index_0[953] = 10'd0;
assign feature_index_0[954] = 10'd0;
assign feature_index_0[955] = 10'd0;
assign feature_index_0[956] = 10'd0;
assign feature_index_0[957] = 10'd597;
assign feature_index_0[958] = 10'd435;
assign feature_index_0[959] = 10'd264;
assign feature_index_0[960] = 10'd159;
assign feature_index_0[961] = 10'd656;
assign feature_index_0[962] = 10'd598;
assign feature_index_0[963] = 10'd706;
assign feature_index_0[964] = 10'd458;
assign feature_index_0[965] = 10'd376;
assign feature_index_0[966] = 10'd513;
assign feature_index_0[967] = 10'd349;
assign feature_index_0[968] = 10'd456;
assign feature_index_0[969] = 10'd434;
assign feature_index_0[970] = 10'd655;
assign feature_index_0[971] = 10'd656;
assign feature_index_0[972] = 10'd598;
assign feature_index_0[973] = 10'd548;
assign feature_index_0[974] = 10'd381;
assign feature_index_0[975] = 10'd210;
assign feature_index_0[976] = 10'd236;
assign feature_index_0[977] = 10'd268;
assign feature_index_0[978] = 10'd298;
assign feature_index_0[979] = 10'd330;
assign feature_index_0[980] = 10'd0;
assign feature_index_0[981] = 10'd0;
assign feature_index_0[982] = 10'd135;
assign feature_index_0[983] = 10'd656;
assign feature_index_0[984] = 10'd524;
assign feature_index_0[985] = 10'd487;
assign feature_index_0[986] = 10'd490;
assign feature_index_0[987] = 10'd347;
assign feature_index_0[988] = 10'd664;
assign feature_index_0[989] = 10'd499;
assign feature_index_0[990] = 10'd512;
assign feature_index_0[991] = 10'd187;
assign feature_index_0[992] = 10'd578;
assign feature_index_0[993] = 10'd379;
assign feature_index_0[994] = 10'd574;
assign feature_index_0[995] = 10'd96;
assign feature_index_0[996] = 10'd576;
assign feature_index_0[997] = 10'd627;
assign feature_index_0[998] = 10'd379;
assign feature_index_0[999] = 10'd181;
assign feature_index_0[1000] = 10'd606;
assign feature_index_0[1001] = 10'd460;
assign feature_index_0[1002] = 10'd372;
assign feature_index_0[1003] = 10'd546;
assign feature_index_0[1004] = 10'd299;
assign feature_index_0[1005] = 10'd233;
assign feature_index_0[1006] = 10'd467;
assign feature_index_0[1007] = 10'd0;
assign feature_index_0[1008] = 10'd0;
assign feature_index_0[1009] = 10'd552;
assign feature_index_0[1010] = 10'd407;
assign feature_index_0[1011] = 10'd464;
assign feature_index_0[1012] = 10'd263;
assign feature_index_0[1013] = 10'd494;
assign feature_index_0[1014] = 10'd260;
assign feature_index_0[1015] = 10'd487;
assign feature_index_0[1016] = 10'd345;
assign feature_index_0[1017] = 10'd158;
assign feature_index_0[1018] = 10'd330;
assign feature_index_0[1019] = 10'd240;
assign feature_index_0[1020] = 10'd603;
assign feature_index_0[1021] = 10'd433;
assign feature_index_0[1022] = 10'd483;
assign feature_index_1[0] = 10'd377;
assign feature_index_1[1] = 10'd153;
assign feature_index_1[2] = 10'd178;
assign feature_index_1[3] = 10'd238;
assign feature_index_1[4] = 10'd409;
assign feature_index_1[5] = 10'd403;
assign feature_index_1[6] = 10'd461;
assign feature_index_1[7] = 10'd465;
assign feature_index_1[8] = 10'd510;
assign feature_index_1[9] = 10'd344;
assign feature_index_1[10] = 10'd598;
assign feature_index_1[11] = 10'd461;
assign feature_index_1[12] = 10'd101;
assign feature_index_1[13] = 10'd291;
assign feature_index_1[14] = 10'd316;
assign feature_index_1[15] = 10'd378;
assign feature_index_1[16] = 10'd295;
assign feature_index_1[17] = 10'd569;
assign feature_index_1[18] = 10'd625;
assign feature_index_1[19] = 10'd271;
assign feature_index_1[20] = 10'd432;
assign feature_index_1[21] = 10'd544;
assign feature_index_1[22] = 10'd412;
assign feature_index_1[23] = 10'd316;
assign feature_index_1[24] = 10'd291;
assign feature_index_1[25] = 10'd488;
assign feature_index_1[26] = 10'd293;
assign feature_index_1[27] = 10'd181;
assign feature_index_1[28] = 10'd176;
assign feature_index_1[29] = 10'd498;
assign feature_index_1[30] = 10'd484;
assign feature_index_1[31] = 10'd323;
assign feature_index_1[32] = 10'd428;
assign feature_index_1[33] = 10'd570;
assign feature_index_1[34] = 10'd293;
assign feature_index_1[35] = 10'd373;
assign feature_index_1[36] = 10'd625;
assign feature_index_1[37] = 10'd381;
assign feature_index_1[38] = 10'd432;
assign feature_index_1[39] = 10'd462;
assign feature_index_1[40] = 10'd461;
assign feature_index_1[41] = 10'd352;
assign feature_index_1[42] = 10'd658;
assign feature_index_1[43] = 10'd681;
assign feature_index_1[44] = 10'd215;
assign feature_index_1[45] = 10'd348;
assign feature_index_1[46] = 10'd272;
assign feature_index_1[47] = 10'd298;
assign feature_index_1[48] = 10'd299;
assign feature_index_1[49] = 10'd329;
assign feature_index_1[50] = 10'd488;
assign feature_index_1[51] = 10'd596;
assign feature_index_1[52] = 10'd327;
assign feature_index_1[53] = 10'd187;
assign feature_index_1[54] = 10'd183;
assign feature_index_1[55] = 10'd233;
assign feature_index_1[56] = 10'd323;
assign feature_index_1[57] = 10'd515;
assign feature_index_1[58] = 10'd513;
assign feature_index_1[59] = 10'd318;
assign feature_index_1[60] = 10'd500;
assign feature_index_1[61] = 10'd544;
assign feature_index_1[62] = 10'd213;
assign feature_index_1[63] = 10'd497;
assign feature_index_1[64] = 10'd568;
assign feature_index_1[65] = 10'd402;
assign feature_index_1[66] = 10'd524;
assign feature_index_1[67] = 10'd429;
assign feature_index_1[68] = 10'd244;
assign feature_index_1[69] = 10'd713;
assign feature_index_1[70] = 10'd151;
assign feature_index_1[71] = 10'd432;
assign feature_index_1[72] = 10'd405;
assign feature_index_1[73] = 10'd234;
assign feature_index_1[74] = 10'd456;
assign feature_index_1[75] = 10'd398;
assign feature_index_1[76] = 10'd412;
assign feature_index_1[77] = 10'd104;
assign feature_index_1[78] = 10'd347;
assign feature_index_1[79] = 10'd217;
assign feature_index_1[80] = 10'd375;
assign feature_index_1[81] = 10'd545;
assign feature_index_1[82] = 10'd349;
assign feature_index_1[83] = 10'd413;
assign feature_index_1[84] = 10'd484;
assign feature_index_1[85] = 10'd357;
assign feature_index_1[86] = 10'd354;
assign feature_index_1[87] = 10'd213;
assign feature_index_1[88] = 10'd513;
assign feature_index_1[89] = 10'd568;
assign feature_index_1[90] = 10'd319;
assign feature_index_1[91] = 10'd289;
assign feature_index_1[92] = 10'd273;
assign feature_index_1[93] = 10'd655;
assign feature_index_1[94] = 10'd655;
assign feature_index_1[95] = 10'd628;
assign feature_index_1[96] = 10'd129;
assign feature_index_1[97] = 10'd380;
assign feature_index_1[98] = 10'd438;
assign feature_index_1[99] = 10'd328;
assign feature_index_1[100] = 10'd441;
assign feature_index_1[101] = 10'd180;
assign feature_index_1[102] = 10'd401;
assign feature_index_1[103] = 10'd519;
assign feature_index_1[104] = 10'd248;
assign feature_index_1[105] = 10'd347;
assign feature_index_1[106] = 10'd212;
assign feature_index_1[107] = 10'd214;
assign feature_index_1[108] = 10'd463;
assign feature_index_1[109] = 10'd628;
assign feature_index_1[110] = 10'd555;
assign feature_index_1[111] = 10'd636;
assign feature_index_1[112] = 10'd542;
assign feature_index_1[113] = 10'd287;
assign feature_index_1[114] = 10'd459;
assign feature_index_1[115] = 10'd270;
assign feature_index_1[116] = 10'd184;
assign feature_index_1[117] = 10'd233;
assign feature_index_1[118] = 10'd164;
assign feature_index_1[119] = 10'd554;
assign feature_index_1[120] = 10'd665;
assign feature_index_1[121] = 10'd483;
assign feature_index_1[122] = 10'd523;
assign feature_index_1[123] = 10'd656;
assign feature_index_1[124] = 10'd69;
assign feature_index_1[125] = 10'd152;
assign feature_index_1[126] = 10'd182;
assign feature_index_1[127] = 10'd128;
assign feature_index_1[128] = 10'd95;
assign feature_index_1[129] = 10'd305;
assign feature_index_1[130] = 10'd374;
assign feature_index_1[131] = 10'd209;
assign feature_index_1[132] = 10'd150;
assign feature_index_1[133] = 10'd329;
assign feature_index_1[134] = 10'd95;
assign feature_index_1[135] = 10'd180;
assign feature_index_1[136] = 10'd184;
assign feature_index_1[137] = 10'd442;
assign feature_index_1[138] = 10'd593;
assign feature_index_1[139] = 10'd429;
assign feature_index_1[140] = 10'd187;
assign feature_index_1[141] = 10'd382;
assign feature_index_1[142] = 10'd178;
assign feature_index_1[143] = 10'd456;
assign feature_index_1[144] = 10'd545;
assign feature_index_1[145] = 10'd401;
assign feature_index_1[146] = 10'd380;
assign feature_index_1[147] = 10'd246;
assign feature_index_1[148] = 10'd465;
assign feature_index_1[149] = 10'd681;
assign feature_index_1[150] = 10'd101;
assign feature_index_1[151] = 10'd320;
assign feature_index_1[152] = 10'd465;
assign feature_index_1[153] = 10'd431;
assign feature_index_1[154] = 10'd262;
assign feature_index_1[155] = 10'd460;
assign feature_index_1[156] = 10'd243;
assign feature_index_1[157] = 10'd456;
assign feature_index_1[158] = 10'd434;
assign feature_index_1[159] = 10'd402;
assign feature_index_1[160] = 10'd656;
assign feature_index_1[161] = 10'd540;
assign feature_index_1[162] = 10'd291;
assign feature_index_1[163] = 10'd595;
assign feature_index_1[164] = 10'd263;
assign feature_index_1[165] = 10'd374;
assign feature_index_1[166] = 10'd263;
assign feature_index_1[167] = 10'd387;
assign feature_index_1[168] = 10'd491;
assign feature_index_1[169] = 10'd273;
assign feature_index_1[170] = 10'd183;
assign feature_index_1[171] = 10'd488;
assign feature_index_1[172] = 10'd464;
assign feature_index_1[173] = 10'd542;
assign feature_index_1[174] = 10'd411;
assign feature_index_1[175] = 10'd318;
assign feature_index_1[176] = 10'd654;
assign feature_index_1[177] = 10'd242;
assign feature_index_1[178] = 10'd176;
assign feature_index_1[179] = 10'd274;
assign feature_index_1[180] = 10'd469;
assign feature_index_1[181] = 10'd316;
assign feature_index_1[182] = 10'd429;
assign feature_index_1[183] = 10'd293;
assign feature_index_1[184] = 10'd683;
assign feature_index_1[185] = 10'd123;
assign feature_index_1[186] = 10'd380;
assign feature_index_1[187] = 10'd269;
assign feature_index_1[188] = 10'd270;
assign feature_index_1[189] = 10'd344;
assign feature_index_1[190] = 10'd461;
assign feature_index_1[191] = 10'd572;
assign feature_index_1[192] = 10'd121;
assign feature_index_1[193] = 10'd181;
assign feature_index_1[194] = 10'd567;
assign feature_index_1[195] = 10'd469;
assign feature_index_1[196] = 10'd294;
assign feature_index_1[197] = 10'd551;
assign feature_index_1[198] = 10'd258;
assign feature_index_1[199] = 10'd262;
assign feature_index_1[200] = 10'd184;
assign feature_index_1[201] = 10'd498;
assign feature_index_1[202] = 10'd371;
assign feature_index_1[203] = 10'd156;
assign feature_index_1[204] = 10'd325;
assign feature_index_1[205] = 10'd156;
assign feature_index_1[206] = 10'd97;
assign feature_index_1[207] = 10'd297;
assign feature_index_1[208] = 10'd570;
assign feature_index_1[209] = 10'd512;
assign feature_index_1[210] = 10'd386;
assign feature_index_1[211] = 10'd526;
assign feature_index_1[212] = 10'd297;
assign feature_index_1[213] = 10'd469;
assign feature_index_1[214] = 10'd434;
assign feature_index_1[215] = 10'd624;
assign feature_index_1[216] = 10'd462;
assign feature_index_1[217] = 10'd467;
assign feature_index_1[218] = 10'd294;
assign feature_index_1[219] = 10'd571;
assign feature_index_1[220] = 10'd455;
assign feature_index_1[221] = 10'd564;
assign feature_index_1[222] = 10'd439;
assign feature_index_1[223] = 10'd630;
assign feature_index_1[224] = 10'd405;
assign feature_index_1[225] = 10'd152;
assign feature_index_1[226] = 10'd663;
assign feature_index_1[227] = 10'd656;
assign feature_index_1[228] = 10'd327;
assign feature_index_1[229] = 10'd692;
assign feature_index_1[230] = 10'd487;
assign feature_index_1[231] = 10'd295;
assign feature_index_1[232] = 10'd653;
assign feature_index_1[233] = 10'd215;
assign feature_index_1[234] = 10'd546;
assign feature_index_1[235] = 10'd292;
assign feature_index_1[236] = 10'd290;
assign feature_index_1[237] = 10'd234;
assign feature_index_1[238] = 10'd0;
assign feature_index_1[239] = 10'd656;
assign feature_index_1[240] = 10'd125;
assign feature_index_1[241] = 10'd95;
assign feature_index_1[242] = 10'd684;
assign feature_index_1[243] = 10'd184;
assign feature_index_1[244] = 10'd606;
assign feature_index_1[245] = 10'd331;
assign feature_index_1[246] = 10'd369;
assign feature_index_1[247] = 10'd455;
assign feature_index_1[248] = 10'd355;
assign feature_index_1[249] = 10'd398;
assign feature_index_1[250] = 10'd0;
assign feature_index_1[251] = 10'd570;
assign feature_index_1[252] = 10'd544;
assign feature_index_1[253] = 10'd313;
assign feature_index_1[254] = 10'd247;
assign feature_index_1[255] = 10'd183;
assign feature_index_1[256] = 10'd490;
assign feature_index_1[257] = 10'd629;
assign feature_index_1[258] = 10'd185;
assign feature_index_1[259] = 10'd294;
assign feature_index_1[260] = 10'd0;
assign feature_index_1[261] = 10'd291;
assign feature_index_1[262] = 10'd441;
assign feature_index_1[263] = 10'd232;
assign feature_index_1[264] = 10'd549;
assign feature_index_1[265] = 10'd300;
assign feature_index_1[266] = 10'd0;
assign feature_index_1[267] = 10'd400;
assign feature_index_1[268] = 10'd659;
assign feature_index_1[269] = 10'd411;
assign feature_index_1[270] = 10'd0;
assign feature_index_1[271] = 10'd489;
assign feature_index_1[272] = 10'd209;
assign feature_index_1[273] = 10'd93;
assign feature_index_1[274] = 10'd186;
assign feature_index_1[275] = 10'd241;
assign feature_index_1[276] = 10'd160;
assign feature_index_1[277] = 10'd290;
assign feature_index_1[278] = 10'd343;
assign feature_index_1[279] = 10'd125;
assign feature_index_1[280] = 10'd96;
assign feature_index_1[281] = 10'd319;
assign feature_index_1[282] = 10'd0;
assign feature_index_1[283] = 10'd260;
assign feature_index_1[284] = 10'd540;
assign feature_index_1[285] = 10'd0;
assign feature_index_1[286] = 10'd660;
assign feature_index_1[287] = 10'd232;
assign feature_index_1[288] = 10'd156;
assign feature_index_1[289] = 10'd376;
assign feature_index_1[290] = 10'd232;
assign feature_index_1[291] = 10'd268;
assign feature_index_1[292] = 10'd435;
assign feature_index_1[293] = 10'd356;
assign feature_index_1[294] = 10'd482;
assign feature_index_1[295] = 10'd242;
assign feature_index_1[296] = 10'd402;
assign feature_index_1[297] = 10'd431;
assign feature_index_1[298] = 10'd372;
assign feature_index_1[299] = 10'd430;
assign feature_index_1[300] = 10'd631;
assign feature_index_1[301] = 10'd516;
assign feature_index_1[302] = 10'd491;
assign feature_index_1[303] = 10'd601;
assign feature_index_1[304] = 10'd412;
assign feature_index_1[305] = 10'd717;
assign feature_index_1[306] = 10'd605;
assign feature_index_1[307] = 10'd374;
assign feature_index_1[308] = 10'd372;
assign feature_index_1[309] = 10'd599;
assign feature_index_1[310] = 10'd242;
assign feature_index_1[311] = 10'd99;
assign feature_index_1[312] = 10'd347;
assign feature_index_1[313] = 10'd302;
assign feature_index_1[314] = 10'd301;
assign feature_index_1[315] = 10'd656;
assign feature_index_1[316] = 10'd314;
assign feature_index_1[317] = 10'd330;
assign feature_index_1[318] = 10'd354;
assign feature_index_1[319] = 10'd640;
assign feature_index_1[320] = 10'd658;
assign feature_index_1[321] = 10'd493;
assign feature_index_1[322] = 10'd284;
assign feature_index_1[323] = 10'd631;
assign feature_index_1[324] = 10'd345;
assign feature_index_1[325] = 10'd319;
assign feature_index_1[326] = 10'd656;
assign feature_index_1[327] = 10'd406;
assign feature_index_1[328] = 10'd434;
assign feature_index_1[329] = 10'd516;
assign feature_index_1[330] = 10'd318;
assign feature_index_1[331] = 10'd347;
assign feature_index_1[332] = 10'd348;
assign feature_index_1[333] = 10'd602;
assign feature_index_1[334] = 10'd653;
assign feature_index_1[335] = 10'd100;
assign feature_index_1[336] = 10'd302;
assign feature_index_1[337] = 10'd117;
assign feature_index_1[338] = 10'd595;
assign feature_index_1[339] = 10'd320;
assign feature_index_1[340] = 10'd183;
assign feature_index_1[341] = 10'd575;
assign feature_index_1[342] = 10'd262;
assign feature_index_1[343] = 10'd233;
assign feature_index_1[344] = 10'd601;
assign feature_index_1[345] = 10'd433;
assign feature_index_1[346] = 10'd598;
assign feature_index_1[347] = 10'd301;
assign feature_index_1[348] = 10'd441;
assign feature_index_1[349] = 10'd0;
assign feature_index_1[350] = 10'd269;
assign feature_index_1[351] = 10'd314;
assign feature_index_1[352] = 10'd436;
assign feature_index_1[353] = 10'd233;
assign feature_index_1[354] = 10'd513;
assign feature_index_1[355] = 10'd235;
assign feature_index_1[356] = 10'd149;
assign feature_index_1[357] = 10'd574;
assign feature_index_1[358] = 10'd0;
assign feature_index_1[359] = 10'd241;
assign feature_index_1[360] = 10'd636;
assign feature_index_1[361] = 10'd322;
assign feature_index_1[362] = 10'd186;
assign feature_index_1[363] = 10'd683;
assign feature_index_1[364] = 10'd634;
assign feature_index_1[365] = 10'd566;
assign feature_index_1[366] = 10'd211;
assign feature_index_1[367] = 10'd290;
assign feature_index_1[368] = 10'd321;
assign feature_index_1[369] = 10'd414;
assign feature_index_1[370] = 10'd432;
assign feature_index_1[371] = 10'd625;
assign feature_index_1[372] = 10'd434;
assign feature_index_1[373] = 10'd404;
assign feature_index_1[374] = 10'd355;
assign feature_index_1[375] = 10'd436;
assign feature_index_1[376] = 10'd345;
assign feature_index_1[377] = 10'd487;
assign feature_index_1[378] = 10'd401;
assign feature_index_1[379] = 10'd629;
assign feature_index_1[380] = 10'd241;
assign feature_index_1[381] = 10'd622;
assign feature_index_1[382] = 10'd373;
assign feature_index_1[383] = 10'd376;
assign feature_index_1[384] = 10'd429;
assign feature_index_1[385] = 10'd122;
assign feature_index_1[386] = 10'd488;
assign feature_index_1[387] = 10'd210;
assign feature_index_1[388] = 10'd653;
assign feature_index_1[389] = 10'd515;
assign feature_index_1[390] = 10'd319;
assign feature_index_1[391] = 10'd435;
assign feature_index_1[392] = 10'd407;
assign feature_index_1[393] = 10'd743;
assign feature_index_1[394] = 10'd159;
assign feature_index_1[395] = 10'd408;
assign feature_index_1[396] = 10'd714;
assign feature_index_1[397] = 10'd314;
assign feature_index_1[398] = 10'd355;
assign feature_index_1[399] = 10'd521;
assign feature_index_1[400] = 10'd208;
assign feature_index_1[401] = 10'd207;
assign feature_index_1[402] = 10'd265;
assign feature_index_1[403] = 10'd381;
assign feature_index_1[404] = 10'd0;
assign feature_index_1[405] = 10'd548;
assign feature_index_1[406] = 10'd594;
assign feature_index_1[407] = 10'd219;
assign feature_index_1[408] = 10'd326;
assign feature_index_1[409] = 10'd567;
assign feature_index_1[410] = 10'd486;
assign feature_index_1[411] = 10'd471;
assign feature_index_1[412] = 10'd564;
assign feature_index_1[413] = 10'd540;
assign feature_index_1[414] = 10'd0;
assign feature_index_1[415] = 10'd687;
assign feature_index_1[416] = 10'd680;
assign feature_index_1[417] = 10'd191;
assign feature_index_1[418] = 10'd654;
assign feature_index_1[419] = 10'd292;
assign feature_index_1[420] = 10'd351;
assign feature_index_1[421] = 10'd241;
assign feature_index_1[422] = 10'd608;
assign feature_index_1[423] = 10'd549;
assign feature_index_1[424] = 10'd285;
assign feature_index_1[425] = 10'd192;
assign feature_index_1[426] = 10'd604;
assign feature_index_1[427] = 10'd438;
assign feature_index_1[428] = 10'd218;
assign feature_index_1[429] = 10'd576;
assign feature_index_1[430] = 10'd628;
assign feature_index_1[431] = 10'd134;
assign feature_index_1[432] = 10'd631;
assign feature_index_1[433] = 10'd623;
assign feature_index_1[434] = 10'd569;
assign feature_index_1[435] = 10'd513;
assign feature_index_1[436] = 10'd353;
assign feature_index_1[437] = 10'd331;
assign feature_index_1[438] = 10'd515;
assign feature_index_1[439] = 10'd157;
assign feature_index_1[440] = 10'd0;
assign feature_index_1[441] = 10'd215;
assign feature_index_1[442] = 10'd399;
assign feature_index_1[443] = 10'd595;
assign feature_index_1[444] = 10'd628;
assign feature_index_1[445] = 10'd0;
assign feature_index_1[446] = 10'd345;
assign feature_index_1[447] = 10'd485;
assign feature_index_1[448] = 10'd259;
assign feature_index_1[449] = 10'd287;
assign feature_index_1[450] = 10'd469;
assign feature_index_1[451] = 10'd598;
assign feature_index_1[452] = 10'd372;
assign feature_index_1[453] = 10'd126;
assign feature_index_1[454] = 10'd603;
assign feature_index_1[455] = 10'd546;
assign feature_index_1[456] = 10'd262;
assign feature_index_1[457] = 10'd492;
assign feature_index_1[458] = 10'd707;
assign feature_index_1[459] = 10'd233;
assign feature_index_1[460] = 10'd414;
assign feature_index_1[461] = 10'd316;
assign feature_index_1[462] = 10'd343;
assign feature_index_1[463] = 10'd490;
assign feature_index_1[464] = 10'd486;
assign feature_index_1[465] = 10'd598;
assign feature_index_1[466] = 10'd323;
assign feature_index_1[467] = 10'd659;
assign feature_index_1[468] = 10'd266;
assign feature_index_1[469] = 10'd237;
assign feature_index_1[470] = 10'd246;
assign feature_index_1[471] = 10'd537;
assign feature_index_1[472] = 10'd542;
assign feature_index_1[473] = 10'd375;
assign feature_index_1[474] = 10'd266;
assign feature_index_1[475] = 10'd599;
assign feature_index_1[476] = 10'd427;
assign feature_index_1[477] = 10'd0;
assign feature_index_1[478] = 10'd0;
assign feature_index_1[479] = 10'd292;
assign feature_index_1[480] = 10'd570;
assign feature_index_1[481] = 10'd438;
assign feature_index_1[482] = 10'd521;
assign feature_index_1[483] = 10'd628;
assign feature_index_1[484] = 10'd0;
assign feature_index_1[485] = 10'd465;
assign feature_index_1[486] = 10'd382;
assign feature_index_1[487] = 10'd660;
assign feature_index_1[488] = 10'd634;
assign feature_index_1[489] = 10'd596;
assign feature_index_1[490] = 10'd489;
assign feature_index_1[491] = 10'd273;
assign feature_index_1[492] = 10'd230;
assign feature_index_1[493] = 10'd681;
assign feature_index_1[494] = 10'd0;
assign feature_index_1[495] = 10'd208;
assign feature_index_1[496] = 10'd209;
assign feature_index_1[497] = 10'd324;
assign feature_index_1[498] = 10'd513;
assign feature_index_1[499] = 10'd179;
assign feature_index_1[500] = 10'd609;
assign feature_index_1[501] = 10'd0;
assign feature_index_1[502] = 10'd0;
assign feature_index_1[503] = 10'd211;
assign feature_index_1[504] = 10'd325;
assign feature_index_1[505] = 10'd123;
assign feature_index_1[506] = 10'd229;
assign feature_index_1[507] = 10'd543;
assign feature_index_1[508] = 10'd273;
assign feature_index_1[509] = 10'd272;
assign feature_index_1[510] = 10'd350;
assign feature_index_1[511] = 10'd205;
assign feature_index_1[512] = 10'd159;
assign feature_index_1[513] = 10'd564;
assign feature_index_1[514] = 10'd259;
assign feature_index_1[515] = 10'd549;
assign feature_index_1[516] = 10'd460;
assign feature_index_1[517] = 10'd631;
assign feature_index_1[518] = 10'd518;
assign feature_index_1[519] = 10'd177;
assign feature_index_1[520] = 10'd289;
assign feature_index_1[521] = 10'd0;
assign feature_index_1[522] = 10'd0;
assign feature_index_1[523] = 10'd442;
assign feature_index_1[524] = 10'd486;
assign feature_index_1[525] = 10'd354;
assign feature_index_1[526] = 10'd382;
assign feature_index_1[527] = 10'd510;
assign feature_index_1[528] = 10'd631;
assign feature_index_1[529] = 10'd246;
assign feature_index_1[530] = 10'd375;
assign feature_index_1[531] = 10'd607;
assign feature_index_1[532] = 10'd734;
assign feature_index_1[533] = 10'd0;
assign feature_index_1[534] = 10'd0;
assign feature_index_1[535] = 10'd571;
assign feature_index_1[536] = 10'd545;
assign feature_index_1[537] = 10'd0;
assign feature_index_1[538] = 10'd0;
assign feature_index_1[539] = 10'd300;
assign feature_index_1[540] = 10'd202;
assign feature_index_1[541] = 10'd0;
assign feature_index_1[542] = 10'd0;
assign feature_index_1[543] = 10'd416;
assign feature_index_1[544] = 10'd359;
assign feature_index_1[545] = 10'd317;
assign feature_index_1[546] = 10'd398;
assign feature_index_1[547] = 10'd90;
assign feature_index_1[548] = 10'd192;
assign feature_index_1[549] = 10'd208;
assign feature_index_1[550] = 10'd600;
assign feature_index_1[551] = 10'd245;
assign feature_index_1[552] = 10'd184;
assign feature_index_1[553] = 10'd149;
assign feature_index_1[554] = 10'd317;
assign feature_index_1[555] = 10'd158;
assign feature_index_1[556] = 10'd429;
assign feature_index_1[557] = 10'd0;
assign feature_index_1[558] = 10'd0;
assign feature_index_1[559] = 10'd352;
assign feature_index_1[560] = 10'd0;
assign feature_index_1[561] = 10'd439;
assign feature_index_1[562] = 10'd433;
assign feature_index_1[563] = 10'd547;
assign feature_index_1[564] = 10'd298;
assign feature_index_1[565] = 10'd0;
assign feature_index_1[566] = 10'd0;
assign feature_index_1[567] = 10'd186;
assign feature_index_1[568] = 10'd403;
assign feature_index_1[569] = 10'd163;
assign feature_index_1[570] = 10'd129;
assign feature_index_1[571] = 10'd0;
assign feature_index_1[572] = 10'd0;
assign feature_index_1[573] = 10'd243;
assign feature_index_1[574] = 10'd0;
assign feature_index_1[575] = 10'd184;
assign feature_index_1[576] = 10'd695;
assign feature_index_1[577] = 10'd555;
assign feature_index_1[578] = 10'd624;
assign feature_index_1[579] = 10'd328;
assign feature_index_1[580] = 10'd571;
assign feature_index_1[581] = 10'd543;
assign feature_index_1[582] = 10'd369;
assign feature_index_1[583] = 10'd398;
assign feature_index_1[584] = 10'd266;
assign feature_index_1[585] = 10'd193;
assign feature_index_1[586] = 10'd740;
assign feature_index_1[587] = 10'd381;
assign feature_index_1[588] = 10'd606;
assign feature_index_1[589] = 10'd159;
assign feature_index_1[590] = 10'd288;
assign feature_index_1[591] = 10'd149;
assign feature_index_1[592] = 10'd433;
assign feature_index_1[593] = 10'd434;
assign feature_index_1[594] = 10'd186;
assign feature_index_1[595] = 10'd492;
assign feature_index_1[596] = 10'd523;
assign feature_index_1[597] = 10'd656;
assign feature_index_1[598] = 10'd552;
assign feature_index_1[599] = 10'd435;
assign feature_index_1[600] = 10'd129;
assign feature_index_1[601] = 10'd155;
assign feature_index_1[602] = 10'd460;
assign feature_index_1[603] = 10'd512;
assign feature_index_1[604] = 10'd240;
assign feature_index_1[605] = 10'd405;
assign feature_index_1[606] = 10'd158;
assign feature_index_1[607] = 10'd423;
assign feature_index_1[608] = 10'd438;
assign feature_index_1[609] = 10'd212;
assign feature_index_1[610] = 10'd497;
assign feature_index_1[611] = 10'd266;
assign feature_index_1[612] = 10'd0;
assign feature_index_1[613] = 10'd414;
assign feature_index_1[614] = 10'd213;
assign feature_index_1[615] = 10'd537;
assign feature_index_1[616] = 10'd358;
assign feature_index_1[617] = 10'd314;
assign feature_index_1[618] = 10'd316;
assign feature_index_1[619] = 10'd595;
assign feature_index_1[620] = 10'd157;
assign feature_index_1[621] = 10'd573;
assign feature_index_1[622] = 10'd343;
assign feature_index_1[623] = 10'd353;
assign feature_index_1[624] = 10'd158;
assign feature_index_1[625] = 10'd519;
assign feature_index_1[626] = 10'd352;
assign feature_index_1[627] = 10'd441;
assign feature_index_1[628] = 10'd380;
assign feature_index_1[629] = 10'd496;
assign feature_index_1[630] = 10'd267;
assign feature_index_1[631] = 10'd706;
assign feature_index_1[632] = 10'd262;
assign feature_index_1[633] = 10'd192;
assign feature_index_1[634] = 10'd291;
assign feature_index_1[635] = 10'd184;
assign feature_index_1[636] = 10'd0;
assign feature_index_1[637] = 10'd428;
assign feature_index_1[638] = 10'd246;
assign feature_index_1[639] = 10'd160;
assign feature_index_1[640] = 10'd0;
assign feature_index_1[641] = 10'd473;
assign feature_index_1[642] = 10'd348;
assign feature_index_1[643] = 10'd125;
assign feature_index_1[644] = 10'd518;
assign feature_index_1[645] = 10'd370;
assign feature_index_1[646] = 10'd0;
assign feature_index_1[647] = 10'd569;
assign feature_index_1[648] = 10'd242;
assign feature_index_1[649] = 10'd371;
assign feature_index_1[650] = 10'd292;
assign feature_index_1[651] = 10'd568;
assign feature_index_1[652] = 10'd349;
assign feature_index_1[653] = 10'd515;
assign feature_index_1[654] = 10'd210;
assign feature_index_1[655] = 10'd160;
assign feature_index_1[656] = 10'd0;
assign feature_index_1[657] = 10'd323;
assign feature_index_1[658] = 10'd432;
assign feature_index_1[659] = 10'd233;
assign feature_index_1[660] = 10'd488;
assign feature_index_1[661] = 10'd396;
assign feature_index_1[662] = 10'd328;
assign feature_index_1[663] = 10'd126;
assign feature_index_1[664] = 10'd575;
assign feature_index_1[665] = 10'd485;
assign feature_index_1[666] = 10'd576;
assign feature_index_1[667] = 10'd0;
assign feature_index_1[668] = 10'd430;
assign feature_index_1[669] = 10'd0;
assign feature_index_1[670] = 10'd0;
assign feature_index_1[671] = 10'd134;
assign feature_index_1[672] = 10'd487;
assign feature_index_1[673] = 10'd121;
assign feature_index_1[674] = 10'd288;
assign feature_index_1[675] = 10'd272;
assign feature_index_1[676] = 10'd0;
assign feature_index_1[677] = 10'd272;
assign feature_index_1[678] = 10'd385;
assign feature_index_1[679] = 10'd636;
assign feature_index_1[680] = 10'd378;
assign feature_index_1[681] = 10'd0;
assign feature_index_1[682] = 10'd0;
assign feature_index_1[683] = 10'd572;
assign feature_index_1[684] = 10'd663;
assign feature_index_1[685] = 10'd660;
assign feature_index_1[686] = 10'd519;
assign feature_index_1[687] = 10'd606;
assign feature_index_1[688] = 10'd0;
assign feature_index_1[689] = 10'd216;
assign feature_index_1[690] = 10'd297;
assign feature_index_1[691] = 10'd0;
assign feature_index_1[692] = 10'd0;
assign feature_index_1[693] = 10'd0;
assign feature_index_1[694] = 10'd601;
assign feature_index_1[695] = 10'd215;
assign feature_index_1[696] = 10'd244;
assign feature_index_1[697] = 10'd260;
assign feature_index_1[698] = 10'd0;
assign feature_index_1[699] = 10'd0;
assign feature_index_1[700] = 10'd0;
assign feature_index_1[701] = 10'd213;
assign feature_index_1[702] = 10'd601;
assign feature_index_1[703] = 10'd187;
assign feature_index_1[704] = 10'd625;
assign feature_index_1[705] = 10'd625;
assign feature_index_1[706] = 10'd263;
assign feature_index_1[707] = 10'd348;
assign feature_index_1[708] = 10'd318;
assign feature_index_1[709] = 10'd380;
assign feature_index_1[710] = 10'd628;
assign feature_index_1[711] = 10'd466;
assign feature_index_1[712] = 10'd462;
assign feature_index_1[713] = 10'd546;
assign feature_index_1[714] = 10'd0;
assign feature_index_1[715] = 10'd0;
assign feature_index_1[716] = 10'd159;
assign feature_index_1[717] = 10'd0;
assign feature_index_1[718] = 10'd0;
assign feature_index_1[719] = 10'd318;
assign feature_index_1[720] = 10'd407;
assign feature_index_1[721] = 10'd290;
assign feature_index_1[722] = 10'd0;
assign feature_index_1[723] = 10'd291;
assign feature_index_1[724] = 10'd240;
assign feature_index_1[725] = 10'd324;
assign feature_index_1[726] = 10'd103;
assign feature_index_1[727] = 10'd412;
assign feature_index_1[728] = 10'd634;
assign feature_index_1[729] = 10'd459;
assign feature_index_1[730] = 10'd403;
assign feature_index_1[731] = 10'd469;
assign feature_index_1[732] = 10'd609;
assign feature_index_1[733] = 10'd518;
assign feature_index_1[734] = 10'd543;
assign feature_index_1[735] = 10'd343;
assign feature_index_1[736] = 10'd347;
assign feature_index_1[737] = 10'd347;
assign feature_index_1[738] = 10'd538;
assign feature_index_1[739] = 10'd597;
assign feature_index_1[740] = 10'd386;
assign feature_index_1[741] = 10'd430;
assign feature_index_1[742] = 10'd328;
assign feature_index_1[743] = 10'd626;
assign feature_index_1[744] = 10'd379;
assign feature_index_1[745] = 10'd239;
assign feature_index_1[746] = 10'd457;
assign feature_index_1[747] = 10'd0;
assign feature_index_1[748] = 10'd0;
assign feature_index_1[749] = 10'd0;
assign feature_index_1[750] = 10'd483;
assign feature_index_1[751] = 10'd151;
assign feature_index_1[752] = 10'd244;
assign feature_index_1[753] = 10'd459;
assign feature_index_1[754] = 10'd593;
assign feature_index_1[755] = 10'd329;
assign feature_index_1[756] = 10'd463;
assign feature_index_1[757] = 10'd541;
assign feature_index_1[758] = 10'd436;
assign feature_index_1[759] = 10'd179;
assign feature_index_1[760] = 10'd319;
assign feature_index_1[761] = 10'd414;
assign feature_index_1[762] = 10'd483;
assign feature_index_1[763] = 10'd462;
assign feature_index_1[764] = 10'd179;
assign feature_index_1[765] = 10'd567;
assign feature_index_1[766] = 10'd231;
assign feature_index_1[767] = 10'd579;
assign feature_index_1[768] = 10'd549;
assign feature_index_1[769] = 10'd233;
assign feature_index_1[770] = 10'd154;
assign feature_index_1[771] = 10'd134;
assign feature_index_1[772] = 10'd239;
assign feature_index_1[773] = 10'd0;
assign feature_index_1[774] = 10'd0;
assign feature_index_1[775] = 10'd540;
assign feature_index_1[776] = 10'd439;
assign feature_index_1[777] = 10'd547;
assign feature_index_1[778] = 10'd595;
assign feature_index_1[779] = 10'd458;
assign feature_index_1[780] = 10'd211;
assign feature_index_1[781] = 10'd495;
assign feature_index_1[782] = 10'd133;
assign feature_index_1[783] = 10'd267;
assign feature_index_1[784] = 10'd125;
assign feature_index_1[785] = 10'd0;
assign feature_index_1[786] = 10'd272;
assign feature_index_1[787] = 10'd626;
assign feature_index_1[788] = 10'd0;
assign feature_index_1[789] = 10'd685;
assign feature_index_1[790] = 10'd331;
assign feature_index_1[791] = 10'd564;
assign feature_index_1[792] = 10'd243;
assign feature_index_1[793] = 10'd0;
assign feature_index_1[794] = 10'd245;
assign feature_index_1[795] = 10'd624;
assign feature_index_1[796] = 10'd650;
assign feature_index_1[797] = 10'd235;
assign feature_index_1[798] = 10'd155;
assign feature_index_1[799] = 10'd580;
assign feature_index_1[800] = 10'd486;
assign feature_index_1[801] = 10'd417;
assign feature_index_1[802] = 10'd542;
assign feature_index_1[803] = 10'd128;
assign feature_index_1[804] = 10'd290;
assign feature_index_1[805] = 10'd99;
assign feature_index_1[806] = 10'd320;
assign feature_index_1[807] = 10'd247;
assign feature_index_1[808] = 10'd536;
assign feature_index_1[809] = 10'd0;
assign feature_index_1[810] = 10'd0;
assign feature_index_1[811] = 10'd522;
assign feature_index_1[812] = 10'd344;
assign feature_index_1[813] = 10'd541;
assign feature_index_1[814] = 10'd0;
assign feature_index_1[815] = 10'd743;
assign feature_index_1[816] = 10'd386;
assign feature_index_1[817] = 10'd214;
assign feature_index_1[818] = 10'd456;
assign feature_index_1[819] = 10'd627;
assign feature_index_1[820] = 10'd155;
assign feature_index_1[821] = 10'd459;
assign feature_index_1[822] = 10'd572;
assign feature_index_1[823] = 10'd487;
assign feature_index_1[824] = 10'd0;
assign feature_index_1[825] = 10'd592;
assign feature_index_1[826] = 10'd656;
assign feature_index_1[827] = 10'd437;
assign feature_index_1[828] = 10'd572;
assign feature_index_1[829] = 10'd0;
assign feature_index_1[830] = 10'd0;
assign feature_index_1[831] = 10'd298;
assign feature_index_1[832] = 10'd184;
assign feature_index_1[833] = 10'd486;
assign feature_index_1[834] = 10'd512;
assign feature_index_1[835] = 10'd152;
assign feature_index_1[836] = 10'd240;
assign feature_index_1[837] = 10'd459;
assign feature_index_1[838] = 10'd603;
assign feature_index_1[839] = 10'd298;
assign feature_index_1[840] = 10'd296;
assign feature_index_1[841] = 10'd356;
assign feature_index_1[842] = 10'd485;
assign feature_index_1[843] = 10'd159;
assign feature_index_1[844] = 10'd218;
assign feature_index_1[845] = 10'd245;
assign feature_index_1[846] = 10'd0;
assign feature_index_1[847] = 10'd465;
assign feature_index_1[848] = 10'd210;
assign feature_index_1[849] = 10'd131;
assign feature_index_1[850] = 10'd554;
assign feature_index_1[851] = 10'd655;
assign feature_index_1[852] = 10'd329;
assign feature_index_1[853] = 10'd541;
assign feature_index_1[854] = 10'd402;
assign feature_index_1[855] = 10'd210;
assign feature_index_1[856] = 10'd184;
assign feature_index_1[857] = 10'd574;
assign feature_index_1[858] = 10'd295;
assign feature_index_1[859] = 10'd592;
assign feature_index_1[860] = 10'd375;
assign feature_index_1[861] = 10'd429;
assign feature_index_1[862] = 10'd438;
assign feature_index_1[863] = 10'd127;
assign feature_index_1[864] = 10'd623;
assign feature_index_1[865] = 10'd550;
assign feature_index_1[866] = 10'd592;
assign feature_index_1[867] = 10'd0;
assign feature_index_1[868] = 10'd0;
assign feature_index_1[869] = 10'd0;
assign feature_index_1[870] = 10'd463;
assign feature_index_1[871] = 10'd541;
assign feature_index_1[872] = 10'd355;
assign feature_index_1[873] = 10'd0;
assign feature_index_1[874] = 10'd272;
assign feature_index_1[875] = 10'd296;
assign feature_index_1[876] = 10'd439;
assign feature_index_1[877] = 10'd0;
assign feature_index_1[878] = 10'd184;
assign feature_index_1[879] = 10'd0;
assign feature_index_1[880] = 10'd0;
assign feature_index_1[881] = 10'd0;
assign feature_index_1[882] = 10'd0;
assign feature_index_1[883] = 10'd0;
assign feature_index_1[884] = 10'd0;
assign feature_index_1[885] = 10'd0;
assign feature_index_1[886] = 10'd0;
assign feature_index_1[887] = 10'd246;
assign feature_index_1[888] = 10'd381;
assign feature_index_1[889] = 10'd301;
assign feature_index_1[890] = 10'd270;
assign feature_index_1[891] = 10'd0;
assign feature_index_1[892] = 10'd0;
assign feature_index_1[893] = 10'd0;
assign feature_index_1[894] = 10'd0;
assign feature_index_1[895] = 10'd350;
assign feature_index_1[896] = 10'd206;
assign feature_index_1[897] = 10'd264;
assign feature_index_1[898] = 10'd519;
assign feature_index_1[899] = 10'd0;
assign feature_index_1[900] = 10'd374;
assign feature_index_1[901] = 10'd287;
assign feature_index_1[902] = 10'd0;
assign feature_index_1[903] = 10'd625;
assign feature_index_1[904] = 10'd265;
assign feature_index_1[905] = 10'd317;
assign feature_index_1[906] = 10'd480;
assign feature_index_1[907] = 10'd0;
assign feature_index_1[908] = 10'd443;
assign feature_index_1[909] = 10'd402;
assign feature_index_1[910] = 10'd0;
assign feature_index_1[911] = 10'd529;
assign feature_index_1[912] = 10'd344;
assign feature_index_1[913] = 10'd546;
assign feature_index_1[914] = 10'd327;
assign feature_index_1[915] = 10'd274;
assign feature_index_1[916] = 10'd325;
assign feature_index_1[917] = 10'd660;
assign feature_index_1[918] = 10'd539;
assign feature_index_1[919] = 10'd290;
assign feature_index_1[920] = 10'd295;
assign feature_index_1[921] = 10'd687;
assign feature_index_1[922] = 10'd0;
assign feature_index_1[923] = 10'd484;
assign feature_index_1[924] = 10'd540;
assign feature_index_1[925] = 10'd688;
assign feature_index_1[926] = 10'd608;
assign feature_index_1[927] = 10'd97;
assign feature_index_1[928] = 10'd431;
assign feature_index_1[929] = 10'd440;
assign feature_index_1[930] = 10'd631;
assign feature_index_1[931] = 10'd212;
assign feature_index_1[932] = 10'd416;
assign feature_index_1[933] = 10'd425;
assign feature_index_1[934] = 10'd264;
assign feature_index_1[935] = 10'd433;
assign feature_index_1[936] = 10'd552;
assign feature_index_1[937] = 10'd0;
assign feature_index_1[938] = 10'd433;
assign feature_index_1[939] = 10'd270;
assign feature_index_1[940] = 10'd374;
assign feature_index_1[941] = 10'd242;
assign feature_index_1[942] = 10'd470;
assign feature_index_1[943] = 10'd0;
assign feature_index_1[944] = 10'd0;
assign feature_index_1[945] = 10'd687;
assign feature_index_1[946] = 10'd528;
assign feature_index_1[947] = 10'd155;
assign feature_index_1[948] = 10'd416;
assign feature_index_1[949] = 10'd271;
assign feature_index_1[950] = 10'd213;
assign feature_index_1[951] = 10'd567;
assign feature_index_1[952] = 10'd353;
assign feature_index_1[953] = 10'd431;
assign feature_index_1[954] = 10'd357;
assign feature_index_1[955] = 10'd0;
assign feature_index_1[956] = 10'd0;
assign feature_index_1[957] = 10'd0;
assign feature_index_1[958] = 10'd0;
assign feature_index_1[959] = 10'd127;
assign feature_index_1[960] = 10'd542;
assign feature_index_1[961] = 10'd523;
assign feature_index_1[962] = 10'd403;
assign feature_index_1[963] = 10'd143;
assign feature_index_1[964] = 10'd350;
assign feature_index_1[965] = 10'd0;
assign feature_index_1[966] = 10'd460;
assign feature_index_1[967] = 10'd154;
assign feature_index_1[968] = 10'd487;
assign feature_index_1[969] = 10'd0;
assign feature_index_1[970] = 10'd0;
assign feature_index_1[971] = 10'd0;
assign feature_index_1[972] = 10'd656;
assign feature_index_1[973] = 10'd0;
assign feature_index_1[974] = 10'd0;
assign feature_index_1[975] = 10'd345;
assign feature_index_1[976] = 10'd350;
assign feature_index_1[977] = 10'd273;
assign feature_index_1[978] = 10'd519;
assign feature_index_1[979] = 10'd291;
assign feature_index_1[980] = 10'd0;
assign feature_index_1[981] = 10'd438;
assign feature_index_1[982] = 10'd315;
assign feature_index_1[983] = 10'd683;
assign feature_index_1[984] = 10'd0;
assign feature_index_1[985] = 10'd0;
assign feature_index_1[986] = 10'd0;
assign feature_index_1[987] = 10'd346;
assign feature_index_1[988] = 10'd0;
assign feature_index_1[989] = 10'd0;
assign feature_index_1[990] = 10'd0;
assign feature_index_1[991] = 10'd382;
assign feature_index_1[992] = 10'd577;
assign feature_index_1[993] = 10'd0;
assign feature_index_1[994] = 10'd665;
assign feature_index_1[995] = 10'd331;
assign feature_index_1[996] = 10'd493;
assign feature_index_1[997] = 10'd551;
assign feature_index_1[998] = 10'd565;
assign feature_index_1[999] = 10'd655;
assign feature_index_1[1000] = 10'd67;
assign feature_index_1[1001] = 10'd486;
assign feature_index_1[1002] = 10'd594;
assign feature_index_1[1003] = 10'd0;
assign feature_index_1[1004] = 10'd0;
assign feature_index_1[1005] = 10'd0;
assign feature_index_1[1006] = 10'd0;
assign feature_index_1[1007] = 10'd466;
assign feature_index_1[1008] = 10'd607;
assign feature_index_1[1009] = 10'd528;
assign feature_index_1[1010] = 10'd0;
assign feature_index_1[1011] = 10'd156;
assign feature_index_1[1012] = 10'd578;
assign feature_index_1[1013] = 10'd622;
assign feature_index_1[1014] = 10'd0;
assign feature_index_1[1015] = 10'd209;
assign feature_index_1[1016] = 10'd0;
assign feature_index_1[1017] = 10'd0;
assign feature_index_1[1018] = 10'd0;
assign feature_index_1[1019] = 10'd557;
assign feature_index_1[1020] = 10'd547;
assign feature_index_1[1021] = 10'd690;
assign feature_index_1[1022] = 10'd463;
assign feature_index_2[0] = 10'd625;
assign feature_index_2[1] = 10'd430;
assign feature_index_2[2] = 10'd380;
assign feature_index_2[3] = 10'd382;
assign feature_index_2[4] = 10'd237;
assign feature_index_2[5] = 10'd491;
assign feature_index_2[6] = 10'd515;
assign feature_index_2[7] = 10'd493;
assign feature_index_2[8] = 10'd404;
assign feature_index_2[9] = 10'd155;
assign feature_index_2[10] = 10'd100;
assign feature_index_2[11] = 10'd301;
assign feature_index_2[12] = 10'd439;
assign feature_index_2[13] = 10'd516;
assign feature_index_2[14] = 10'd347;
assign feature_index_2[15] = 10'd406;
assign feature_index_2[16] = 10'd406;
assign feature_index_2[17] = 10'd399;
assign feature_index_2[18] = 10'd237;
assign feature_index_2[19] = 10'd514;
assign feature_index_2[20] = 10'd345;
assign feature_index_2[21] = 10'd571;
assign feature_index_2[22] = 10'd508;
assign feature_index_2[23] = 10'd426;
assign feature_index_2[24] = 10'd236;
assign feature_index_2[25] = 10'd381;
assign feature_index_2[26] = 10'd346;
assign feature_index_2[27] = 10'd511;
assign feature_index_2[28] = 10'd710;
assign feature_index_2[29] = 10'd603;
assign feature_index_2[30] = 10'd440;
assign feature_index_2[31] = 10'd569;
assign feature_index_2[32] = 10'd409;
assign feature_index_2[33] = 10'd274;
assign feature_index_2[34] = 10'd494;
assign feature_index_2[35] = 10'd568;
assign feature_index_2[36] = 10'd524;
assign feature_index_2[37] = 10'd544;
assign feature_index_2[38] = 10'd491;
assign feature_index_2[39] = 10'd567;
assign feature_index_2[40] = 10'd215;
assign feature_index_2[41] = 10'd538;
assign feature_index_2[42] = 10'd627;
assign feature_index_2[43] = 10'd348;
assign feature_index_2[44] = 10'd659;
assign feature_index_2[45] = 10'd214;
assign feature_index_2[46] = 10'd0;
assign feature_index_2[47] = 10'd484;
assign feature_index_2[48] = 10'd433;
assign feature_index_2[49] = 10'd461;
assign feature_index_2[50] = 10'd487;
assign feature_index_2[51] = 10'd351;
assign feature_index_2[52] = 10'd267;
assign feature_index_2[53] = 10'd150;
assign feature_index_2[54] = 10'd511;
assign feature_index_2[55] = 10'd290;
assign feature_index_2[56] = 10'd298;
assign feature_index_2[57] = 10'd512;
assign feature_index_2[58] = 10'd433;
assign feature_index_2[59] = 10'd153;
assign feature_index_2[60] = 10'd581;
assign feature_index_2[61] = 10'd432;
assign feature_index_2[62] = 10'd182;
assign feature_index_2[63] = 10'd377;
assign feature_index_2[64] = 10'd398;
assign feature_index_2[65] = 10'd290;
assign feature_index_2[66] = 10'd405;
assign feature_index_2[67] = 10'd129;
assign feature_index_2[68] = 10'd215;
assign feature_index_2[69] = 10'd125;
assign feature_index_2[70] = 10'd662;
assign feature_index_2[71] = 10'd513;
assign feature_index_2[72] = 10'd461;
assign feature_index_2[73] = 10'd682;
assign feature_index_2[74] = 10'd269;
assign feature_index_2[75] = 10'd492;
assign feature_index_2[76] = 10'd429;
assign feature_index_2[77] = 10'd658;
assign feature_index_2[78] = 10'd433;
assign feature_index_2[79] = 10'd353;
assign feature_index_2[80] = 10'd484;
assign feature_index_2[81] = 10'd576;
assign feature_index_2[82] = 10'd267;
assign feature_index_2[83] = 10'd658;
assign feature_index_2[84] = 10'd604;
assign feature_index_2[85] = 10'd178;
assign feature_index_2[86] = 10'd405;
assign feature_index_2[87] = 10'd241;
assign feature_index_2[88] = 10'd267;
assign feature_index_2[89] = 10'd129;
assign feature_index_2[90] = 10'd513;
assign feature_index_2[91] = 10'd573;
assign feature_index_2[92] = 10'd319;
assign feature_index_2[93] = 10'd0;
assign feature_index_2[94] = 10'd0;
assign feature_index_2[95] = 10'd488;
assign feature_index_2[96] = 10'd456;
assign feature_index_2[97] = 10'd556;
assign feature_index_2[98] = 10'd149;
assign feature_index_2[99] = 10'd524;
assign feature_index_2[100] = 10'd357;
assign feature_index_2[101] = 10'd399;
assign feature_index_2[102] = 10'd186;
assign feature_index_2[103] = 10'd150;
assign feature_index_2[104] = 10'd292;
assign feature_index_2[105] = 10'd329;
assign feature_index_2[106] = 10'd521;
assign feature_index_2[107] = 10'd153;
assign feature_index_2[108] = 10'd347;
assign feature_index_2[109] = 10'd432;
assign feature_index_2[110] = 10'd435;
assign feature_index_2[111] = 10'd550;
assign feature_index_2[112] = 10'd491;
assign feature_index_2[113] = 10'd356;
assign feature_index_2[114] = 10'd484;
assign feature_index_2[115] = 10'd401;
assign feature_index_2[116] = 10'd237;
assign feature_index_2[117] = 10'd240;
assign feature_index_2[118] = 10'd185;
assign feature_index_2[119] = 10'd410;
assign feature_index_2[120] = 10'd345;
assign feature_index_2[121] = 10'd125;
assign feature_index_2[122] = 10'd369;
assign feature_index_2[123] = 10'd378;
assign feature_index_2[124] = 10'd183;
assign feature_index_2[125] = 10'd211;
assign feature_index_2[126] = 10'd460;
assign feature_index_2[127] = 10'd381;
assign feature_index_2[128] = 10'd379;
assign feature_index_2[129] = 10'd320;
assign feature_index_2[130] = 10'd465;
assign feature_index_2[131] = 10'd580;
assign feature_index_2[132] = 10'd551;
assign feature_index_2[133] = 10'd577;
assign feature_index_2[134] = 10'd462;
assign feature_index_2[135] = 10'd375;
assign feature_index_2[136] = 10'd300;
assign feature_index_2[137] = 10'd297;
assign feature_index_2[138] = 10'd441;
assign feature_index_2[139] = 10'd571;
assign feature_index_2[140] = 10'd237;
assign feature_index_2[141] = 10'd489;
assign feature_index_2[142] = 10'd516;
assign feature_index_2[143] = 10'd152;
assign feature_index_2[144] = 10'd345;
assign feature_index_2[145] = 10'd125;
assign feature_index_2[146] = 10'd711;
assign feature_index_2[147] = 10'd487;
assign feature_index_2[148] = 10'd514;
assign feature_index_2[149] = 10'd601;
assign feature_index_2[150] = 10'd515;
assign feature_index_2[151] = 10'd318;
assign feature_index_2[152] = 10'd568;
assign feature_index_2[153] = 10'd631;
assign feature_index_2[154] = 10'd316;
assign feature_index_2[155] = 10'd433;
assign feature_index_2[156] = 10'd434;
assign feature_index_2[157] = 10'd544;
assign feature_index_2[158] = 10'd514;
assign feature_index_2[159] = 10'd320;
assign feature_index_2[160] = 10'd439;
assign feature_index_2[161] = 10'd468;
assign feature_index_2[162] = 10'd349;
assign feature_index_2[163] = 10'd276;
assign feature_index_2[164] = 10'd689;
assign feature_index_2[165] = 10'd596;
assign feature_index_2[166] = 10'd160;
assign feature_index_2[167] = 10'd342;
assign feature_index_2[168] = 10'd263;
assign feature_index_2[169] = 10'd542;
assign feature_index_2[170] = 10'd545;
assign feature_index_2[171] = 10'd181;
assign feature_index_2[172] = 10'd97;
assign feature_index_2[173] = 10'd376;
assign feature_index_2[174] = 10'd327;
assign feature_index_2[175] = 10'd211;
assign feature_index_2[176] = 10'd189;
assign feature_index_2[177] = 10'd325;
assign feature_index_2[178] = 10'd229;
assign feature_index_2[179] = 10'd99;
assign feature_index_2[180] = 10'd273;
assign feature_index_2[181] = 10'd461;
assign feature_index_2[182] = 10'd404;
assign feature_index_2[183] = 10'd541;
assign feature_index_2[184] = 10'd203;
assign feature_index_2[185] = 10'd581;
assign feature_index_2[186] = 10'd300;
assign feature_index_2[187] = 10'd0;
assign feature_index_2[188] = 10'd0;
assign feature_index_2[189] = 10'd0;
assign feature_index_2[190] = 10'd0;
assign feature_index_2[191] = 10'd288;
assign feature_index_2[192] = 10'd434;
assign feature_index_2[193] = 10'd175;
assign feature_index_2[194] = 10'd328;
assign feature_index_2[195] = 10'd248;
assign feature_index_2[196] = 10'd229;
assign feature_index_2[197] = 10'd482;
assign feature_index_2[198] = 10'd327;
assign feature_index_2[199] = 10'd517;
assign feature_index_2[200] = 10'd546;
assign feature_index_2[201] = 10'd231;
assign feature_index_2[202] = 10'd294;
assign feature_index_2[203] = 10'd406;
assign feature_index_2[204] = 10'd461;
assign feature_index_2[205] = 10'd460;
assign feature_index_2[206] = 10'd540;
assign feature_index_2[207] = 10'd104;
assign feature_index_2[208] = 10'd160;
assign feature_index_2[209] = 10'd516;
assign feature_index_2[210] = 10'd154;
assign feature_index_2[211] = 10'd579;
assign feature_index_2[212] = 10'd432;
assign feature_index_2[213] = 10'd461;
assign feature_index_2[214] = 10'd188;
assign feature_index_2[215] = 10'd680;
assign feature_index_2[216] = 10'd351;
assign feature_index_2[217] = 10'd648;
assign feature_index_2[218] = 10'd157;
assign feature_index_2[219] = 10'd288;
assign feature_index_2[220] = 10'd495;
assign feature_index_2[221] = 10'd582;
assign feature_index_2[222] = 10'd298;
assign feature_index_2[223] = 10'd181;
assign feature_index_2[224] = 10'd486;
assign feature_index_2[225] = 10'd345;
assign feature_index_2[226] = 10'd345;
assign feature_index_2[227] = 10'd216;
assign feature_index_2[228] = 10'd431;
assign feature_index_2[229] = 10'd221;
assign feature_index_2[230] = 10'd96;
assign feature_index_2[231] = 10'd603;
assign feature_index_2[232] = 10'd549;
assign feature_index_2[233] = 10'd371;
assign feature_index_2[234] = 10'd245;
assign feature_index_2[235] = 10'd213;
assign feature_index_2[236] = 10'd500;
assign feature_index_2[237] = 10'd267;
assign feature_index_2[238] = 10'd219;
assign feature_index_2[239] = 10'd710;
assign feature_index_2[240] = 10'd594;
assign feature_index_2[241] = 10'd483;
assign feature_index_2[242] = 10'd621;
assign feature_index_2[243] = 10'd635;
assign feature_index_2[244] = 10'd320;
assign feature_index_2[245] = 10'd461;
assign feature_index_2[246] = 10'd435;
assign feature_index_2[247] = 10'd271;
assign feature_index_2[248] = 10'd629;
assign feature_index_2[249] = 10'd104;
assign feature_index_2[250] = 10'd630;
assign feature_index_2[251] = 10'd433;
assign feature_index_2[252] = 10'd131;
assign feature_index_2[253] = 10'd376;
assign feature_index_2[254] = 10'd102;
assign feature_index_2[255] = 10'd296;
assign feature_index_2[256] = 10'd485;
assign feature_index_2[257] = 10'd489;
assign feature_index_2[258] = 10'd435;
assign feature_index_2[259] = 10'd325;
assign feature_index_2[260] = 10'd487;
assign feature_index_2[261] = 10'd599;
assign feature_index_2[262] = 10'd0;
assign feature_index_2[263] = 10'd514;
assign feature_index_2[264] = 10'd454;
assign feature_index_2[265] = 10'd576;
assign feature_index_2[266] = 10'd371;
assign feature_index_2[267] = 10'd462;
assign feature_index_2[268] = 10'd374;
assign feature_index_2[269] = 10'd572;
assign feature_index_2[270] = 10'd260;
assign feature_index_2[271] = 10'd514;
assign feature_index_2[272] = 10'd328;
assign feature_index_2[273] = 10'd269;
assign feature_index_2[274] = 10'd0;
assign feature_index_2[275] = 10'd489;
assign feature_index_2[276] = 10'd467;
assign feature_index_2[277] = 10'd487;
assign feature_index_2[278] = 10'd415;
assign feature_index_2[279] = 10'd353;
assign feature_index_2[280] = 10'd684;
assign feature_index_2[281] = 10'd176;
assign feature_index_2[282] = 10'd295;
assign feature_index_2[283] = 10'd322;
assign feature_index_2[284] = 10'd375;
assign feature_index_2[285] = 10'd261;
assign feature_index_2[286] = 10'd376;
assign feature_index_2[287] = 10'd377;
assign feature_index_2[288] = 10'd348;
assign feature_index_2[289] = 10'd233;
assign feature_index_2[290] = 10'd412;
assign feature_index_2[291] = 10'd329;
assign feature_index_2[292] = 10'd320;
assign feature_index_2[293] = 10'd292;
assign feature_index_2[294] = 10'd546;
assign feature_index_2[295] = 10'd541;
assign feature_index_2[296] = 10'd267;
assign feature_index_2[297] = 10'd688;
assign feature_index_2[298] = 10'd213;
assign feature_index_2[299] = 10'd607;
assign feature_index_2[300] = 10'd609;
assign feature_index_2[301] = 10'd235;
assign feature_index_2[302] = 10'd183;
assign feature_index_2[303] = 10'd692;
assign feature_index_2[304] = 10'd270;
assign feature_index_2[305] = 10'd598;
assign feature_index_2[306] = 10'd514;
assign feature_index_2[307] = 10'd634;
assign feature_index_2[308] = 10'd569;
assign feature_index_2[309] = 10'd629;
assign feature_index_2[310] = 10'd0;
assign feature_index_2[311] = 10'd599;
assign feature_index_2[312] = 10'd493;
assign feature_index_2[313] = 10'd547;
assign feature_index_2[314] = 10'd274;
assign feature_index_2[315] = 10'd541;
assign feature_index_2[316] = 10'd212;
assign feature_index_2[317] = 10'd415;
assign feature_index_2[318] = 10'd583;
assign feature_index_2[319] = 10'd683;
assign feature_index_2[320] = 10'd181;
assign feature_index_2[321] = 10'd207;
assign feature_index_2[322] = 10'd97;
assign feature_index_2[323] = 10'd127;
assign feature_index_2[324] = 10'd0;
assign feature_index_2[325] = 10'd491;
assign feature_index_2[326] = 10'd462;
assign feature_index_2[327] = 10'd104;
assign feature_index_2[328] = 10'd298;
assign feature_index_2[329] = 10'd189;
assign feature_index_2[330] = 10'd374;
assign feature_index_2[331] = 10'd598;
assign feature_index_2[332] = 10'd323;
assign feature_index_2[333] = 10'd158;
assign feature_index_2[334] = 10'd244;
assign feature_index_2[335] = 10'd74;
assign feature_index_2[336] = 10'd516;
assign feature_index_2[337] = 10'd316;
assign feature_index_2[338] = 10'd378;
assign feature_index_2[339] = 10'd628;
assign feature_index_2[340] = 10'd0;
assign feature_index_2[341] = 10'd516;
assign feature_index_2[342] = 10'd244;
assign feature_index_2[343] = 10'd243;
assign feature_index_2[344] = 10'd262;
assign feature_index_2[345] = 10'd576;
assign feature_index_2[346] = 10'd514;
assign feature_index_2[347] = 10'd434;
assign feature_index_2[348] = 10'd455;
assign feature_index_2[349] = 10'd270;
assign feature_index_2[350] = 10'd456;
assign feature_index_2[351] = 10'd272;
assign feature_index_2[352] = 10'd410;
assign feature_index_2[353] = 10'd442;
assign feature_index_2[354] = 10'd272;
assign feature_index_2[355] = 10'd463;
assign feature_index_2[356] = 10'd239;
assign feature_index_2[357] = 10'd271;
assign feature_index_2[358] = 10'd520;
assign feature_index_2[359] = 10'd542;
assign feature_index_2[360] = 10'd243;
assign feature_index_2[361] = 10'd102;
assign feature_index_2[362] = 10'd510;
assign feature_index_2[363] = 10'd635;
assign feature_index_2[364] = 10'd327;
assign feature_index_2[365] = 10'd433;
assign feature_index_2[366] = 10'd407;
assign feature_index_2[367] = 10'd261;
assign feature_index_2[368] = 10'd296;
assign feature_index_2[369] = 10'd557;
assign feature_index_2[370] = 10'd256;
assign feature_index_2[371] = 10'd353;
assign feature_index_2[372] = 10'd0;
assign feature_index_2[373] = 10'd153;
assign feature_index_2[374] = 10'd404;
assign feature_index_2[375] = 10'd0;
assign feature_index_2[376] = 10'd0;
assign feature_index_2[377] = 10'd0;
assign feature_index_2[378] = 10'd0;
assign feature_index_2[379] = 10'd0;
assign feature_index_2[380] = 10'd0;
assign feature_index_2[381] = 10'd0;
assign feature_index_2[382] = 10'd0;
assign feature_index_2[383] = 10'd291;
assign feature_index_2[384] = 10'd474;
assign feature_index_2[385] = 10'd154;
assign feature_index_2[386] = 10'd205;
assign feature_index_2[387] = 10'd100;
assign feature_index_2[388] = 10'd515;
assign feature_index_2[389] = 10'd653;
assign feature_index_2[390] = 10'd405;
assign feature_index_2[391] = 10'd454;
assign feature_index_2[392] = 10'd714;
assign feature_index_2[393] = 10'd0;
assign feature_index_2[394] = 10'd0;
assign feature_index_2[395] = 10'd180;
assign feature_index_2[396] = 10'd318;
assign feature_index_2[397] = 10'd0;
assign feature_index_2[398] = 10'd0;
assign feature_index_2[399] = 10'd406;
assign feature_index_2[400] = 10'd578;
assign feature_index_2[401] = 10'd350;
assign feature_index_2[402] = 10'd212;
assign feature_index_2[403] = 10'd411;
assign feature_index_2[404] = 10'd0;
assign feature_index_2[405] = 10'd158;
assign feature_index_2[406] = 10'd511;
assign feature_index_2[407] = 10'd198;
assign feature_index_2[408] = 10'd413;
assign feature_index_2[409] = 10'd210;
assign feature_index_2[410] = 10'd494;
assign feature_index_2[411] = 10'd546;
assign feature_index_2[412] = 10'd434;
assign feature_index_2[413] = 10'd629;
assign feature_index_2[414] = 10'd320;
assign feature_index_2[415] = 10'd433;
assign feature_index_2[416] = 10'd542;
assign feature_index_2[417] = 10'd545;
assign feature_index_2[418] = 10'd412;
assign feature_index_2[419] = 10'd577;
assign feature_index_2[420] = 10'd601;
assign feature_index_2[421] = 10'd573;
assign feature_index_2[422] = 10'd495;
assign feature_index_2[423] = 10'd289;
assign feature_index_2[424] = 10'd658;
assign feature_index_2[425] = 10'd522;
assign feature_index_2[426] = 10'd302;
assign feature_index_2[427] = 10'd603;
assign feature_index_2[428] = 10'd678;
assign feature_index_2[429] = 10'd543;
assign feature_index_2[430] = 10'd538;
assign feature_index_2[431] = 10'd348;
assign feature_index_2[432] = 10'd461;
assign feature_index_2[433] = 10'd272;
assign feature_index_2[434] = 10'd378;
assign feature_index_2[435] = 10'd690;
assign feature_index_2[436] = 10'd128;
assign feature_index_2[437] = 10'd0;
assign feature_index_2[438] = 10'd0;
assign feature_index_2[439] = 10'd435;
assign feature_index_2[440] = 10'd514;
assign feature_index_2[441] = 10'd456;
assign feature_index_2[442] = 10'd434;
assign feature_index_2[443] = 10'd446;
assign feature_index_2[444] = 10'd436;
assign feature_index_2[445] = 10'd355;
assign feature_index_2[446] = 10'd402;
assign feature_index_2[447] = 10'd126;
assign feature_index_2[448] = 10'd399;
assign feature_index_2[449] = 10'd323;
assign feature_index_2[450] = 10'd206;
assign feature_index_2[451] = 10'd297;
assign feature_index_2[452] = 10'd324;
assign feature_index_2[453] = 10'd432;
assign feature_index_2[454] = 10'd595;
assign feature_index_2[455] = 10'd457;
assign feature_index_2[456] = 10'd104;
assign feature_index_2[457] = 10'd152;
assign feature_index_2[458] = 10'd104;
assign feature_index_2[459] = 10'd381;
assign feature_index_2[460] = 10'd0;
assign feature_index_2[461] = 10'd378;
assign feature_index_2[462] = 10'd343;
assign feature_index_2[463] = 10'd150;
assign feature_index_2[464] = 10'd370;
assign feature_index_2[465] = 10'd212;
assign feature_index_2[466] = 10'd397;
assign feature_index_2[467] = 10'd265;
assign feature_index_2[468] = 10'd216;
assign feature_index_2[469] = 10'd373;
assign feature_index_2[470] = 10'd494;
assign feature_index_2[471] = 10'd325;
assign feature_index_2[472] = 10'd346;
assign feature_index_2[473] = 10'd352;
assign feature_index_2[474] = 10'd0;
assign feature_index_2[475] = 10'd211;
assign feature_index_2[476] = 10'd404;
assign feature_index_2[477] = 10'd377;
assign feature_index_2[478] = 10'd376;
assign feature_index_2[479] = 10'd237;
assign feature_index_2[480] = 10'd269;
assign feature_index_2[481] = 10'd709;
assign feature_index_2[482] = 10'd654;
assign feature_index_2[483] = 10'd548;
assign feature_index_2[484] = 10'd0;
assign feature_index_2[485] = 10'd658;
assign feature_index_2[486] = 10'd0;
assign feature_index_2[487] = 10'd656;
assign feature_index_2[488] = 10'd353;
assign feature_index_2[489] = 10'd345;
assign feature_index_2[490] = 10'd433;
assign feature_index_2[491] = 10'd495;
assign feature_index_2[492] = 10'd403;
assign feature_index_2[493] = 10'd0;
assign feature_index_2[494] = 10'd656;
assign feature_index_2[495] = 10'd494;
assign feature_index_2[496] = 10'd513;
assign feature_index_2[497] = 10'd652;
assign feature_index_2[498] = 10'd490;
assign feature_index_2[499] = 10'd241;
assign feature_index_2[500] = 10'd0;
assign feature_index_2[501] = 10'd456;
assign feature_index_2[502] = 10'd318;
assign feature_index_2[503] = 10'd399;
assign feature_index_2[504] = 10'd487;
assign feature_index_2[505] = 10'd733;
assign feature_index_2[506] = 10'd545;
assign feature_index_2[507] = 10'd128;
assign feature_index_2[508] = 10'd290;
assign feature_index_2[509] = 10'd659;
assign feature_index_2[510] = 10'd374;
assign feature_index_2[511] = 10'd594;
assign feature_index_2[512] = 10'd628;
assign feature_index_2[513] = 10'd578;
assign feature_index_2[514] = 10'd345;
assign feature_index_2[515] = 10'd598;
assign feature_index_2[516] = 10'd552;
assign feature_index_2[517] = 10'd544;
assign feature_index_2[518] = 10'd179;
assign feature_index_2[519] = 10'd410;
assign feature_index_2[520] = 10'd381;
assign feature_index_2[521] = 10'd359;
assign feature_index_2[522] = 10'd103;
assign feature_index_2[523] = 10'd350;
assign feature_index_2[524] = 10'd436;
assign feature_index_2[525] = 10'd0;
assign feature_index_2[526] = 10'd0;
assign feature_index_2[527] = 10'd512;
assign feature_index_2[528] = 10'd273;
assign feature_index_2[529] = 10'd414;
assign feature_index_2[530] = 10'd719;
assign feature_index_2[531] = 10'd517;
assign feature_index_2[532] = 10'd267;
assign feature_index_2[533] = 10'd385;
assign feature_index_2[534] = 10'd264;
assign feature_index_2[535] = 10'd482;
assign feature_index_2[536] = 10'd635;
assign feature_index_2[537] = 10'd688;
assign feature_index_2[538] = 10'd381;
assign feature_index_2[539] = 10'd182;
assign feature_index_2[540] = 10'd439;
assign feature_index_2[541] = 10'd317;
assign feature_index_2[542] = 10'd714;
assign feature_index_2[543] = 10'd598;
assign feature_index_2[544] = 10'd359;
assign feature_index_2[545] = 10'd352;
assign feature_index_2[546] = 10'd569;
assign feature_index_2[547] = 10'd515;
assign feature_index_2[548] = 10'd428;
assign feature_index_2[549] = 10'd0;
assign feature_index_2[550] = 10'd0;
assign feature_index_2[551] = 10'd302;
assign feature_index_2[552] = 10'd129;
assign feature_index_2[553] = 10'd133;
assign feature_index_2[554] = 10'd341;
assign feature_index_2[555] = 10'd568;
assign feature_index_2[556] = 10'd598;
assign feature_index_2[557] = 10'd372;
assign feature_index_2[558] = 10'd541;
assign feature_index_2[559] = 10'd123;
assign feature_index_2[560] = 10'd656;
assign feature_index_2[561] = 10'd181;
assign feature_index_2[562] = 10'd516;
assign feature_index_2[563] = 10'd208;
assign feature_index_2[564] = 10'd0;
assign feature_index_2[565] = 10'd487;
assign feature_index_2[566] = 10'd539;
assign feature_index_2[567] = 10'd327;
assign feature_index_2[568] = 10'd219;
assign feature_index_2[569] = 10'd605;
assign feature_index_2[570] = 10'd428;
assign feature_index_2[571] = 10'd343;
assign feature_index_2[572] = 10'd186;
assign feature_index_2[573] = 10'd550;
assign feature_index_2[574] = 10'd117;
assign feature_index_2[575] = 10'd428;
assign feature_index_2[576] = 10'd257;
assign feature_index_2[577] = 10'd683;
assign feature_index_2[578] = 10'd146;
assign feature_index_2[579] = 10'd491;
assign feature_index_2[580] = 10'd518;
assign feature_index_2[581] = 10'd98;
assign feature_index_2[582] = 10'd496;
assign feature_index_2[583] = 10'd151;
assign feature_index_2[584] = 10'd370;
assign feature_index_2[585] = 10'd519;
assign feature_index_2[586] = 10'd124;
assign feature_index_2[587] = 10'd464;
assign feature_index_2[588] = 10'd401;
assign feature_index_2[589] = 10'd0;
assign feature_index_2[590] = 10'd0;
assign feature_index_2[591] = 10'd548;
assign feature_index_2[592] = 10'd214;
assign feature_index_2[593] = 10'd247;
assign feature_index_2[594] = 10'd236;
assign feature_index_2[595] = 10'd221;
assign feature_index_2[596] = 10'd599;
assign feature_index_2[597] = 10'd0;
assign feature_index_2[598] = 10'd628;
assign feature_index_2[599] = 10'd549;
assign feature_index_2[600] = 10'd323;
assign feature_index_2[601] = 10'd551;
assign feature_index_2[602] = 10'd455;
assign feature_index_2[603] = 10'd379;
assign feature_index_2[604] = 10'd656;
assign feature_index_2[605] = 10'd456;
assign feature_index_2[606] = 10'd411;
assign feature_index_2[607] = 10'd657;
assign feature_index_2[608] = 10'd584;
assign feature_index_2[609] = 10'd488;
assign feature_index_2[610] = 10'd208;
assign feature_index_2[611] = 10'd497;
assign feature_index_2[612] = 10'd656;
assign feature_index_2[613] = 10'd177;
assign feature_index_2[614] = 10'd0;
assign feature_index_2[615] = 10'd656;
assign feature_index_2[616] = 10'd688;
assign feature_index_2[617] = 10'd157;
assign feature_index_2[618] = 10'd300;
assign feature_index_2[619] = 10'd0;
assign feature_index_2[620] = 10'd411;
assign feature_index_2[621] = 10'd0;
assign feature_index_2[622] = 10'd0;
assign feature_index_2[623] = 10'd316;
assign feature_index_2[624] = 10'd580;
assign feature_index_2[625] = 10'd400;
assign feature_index_2[626] = 10'd322;
assign feature_index_2[627] = 10'd158;
assign feature_index_2[628] = 10'd379;
assign feature_index_2[629] = 10'd571;
assign feature_index_2[630] = 10'd517;
assign feature_index_2[631] = 10'd689;
assign feature_index_2[632] = 10'd0;
assign feature_index_2[633] = 10'd463;
assign feature_index_2[634] = 10'd601;
assign feature_index_2[635] = 10'd178;
assign feature_index_2[636] = 10'd129;
assign feature_index_2[637] = 10'd657;
assign feature_index_2[638] = 10'd443;
assign feature_index_2[639] = 10'd94;
assign feature_index_2[640] = 10'd384;
assign feature_index_2[641] = 10'd296;
assign feature_index_2[642] = 10'd98;
assign feature_index_2[643] = 10'd266;
assign feature_index_2[644] = 10'd178;
assign feature_index_2[645] = 10'd741;
assign feature_index_2[646] = 10'd0;
assign feature_index_2[647] = 10'd295;
assign feature_index_2[648] = 10'd0;
assign feature_index_2[649] = 10'd0;
assign feature_index_2[650] = 10'd0;
assign feature_index_2[651] = 10'd603;
assign feature_index_2[652] = 10'd464;
assign feature_index_2[653] = 10'd412;
assign feature_index_2[654] = 10'd158;
assign feature_index_2[655] = 10'd437;
assign feature_index_2[656] = 10'd270;
assign feature_index_2[657] = 10'd325;
assign feature_index_2[658] = 10'd469;
assign feature_index_2[659] = 10'd688;
assign feature_index_2[660] = 10'd463;
assign feature_index_2[661] = 10'd207;
assign feature_index_2[662] = 10'd634;
assign feature_index_2[663] = 10'd239;
assign feature_index_2[664] = 10'd353;
assign feature_index_2[665] = 10'd207;
assign feature_index_2[666] = 10'd572;
assign feature_index_2[667] = 10'd386;
assign feature_index_2[668] = 10'd600;
assign feature_index_2[669] = 10'd350;
assign feature_index_2[670] = 10'd352;
assign feature_index_2[671] = 10'd97;
assign feature_index_2[672] = 10'd0;
assign feature_index_2[673] = 10'd269;
assign feature_index_2[674] = 10'd443;
assign feature_index_2[675] = 10'd543;
assign feature_index_2[676] = 10'd288;
assign feature_index_2[677] = 10'd291;
assign feature_index_2[678] = 10'd349;
assign feature_index_2[679] = 10'd0;
assign feature_index_2[680] = 10'd0;
assign feature_index_2[681] = 10'd0;
assign feature_index_2[682] = 10'd0;
assign feature_index_2[683] = 10'd0;
assign feature_index_2[684] = 10'd0;
assign feature_index_2[685] = 10'd466;
assign feature_index_2[686] = 10'd0;
assign feature_index_2[687] = 10'd95;
assign feature_index_2[688] = 10'd538;
assign feature_index_2[689] = 10'd657;
assign feature_index_2[690] = 10'd440;
assign feature_index_2[691] = 10'd469;
assign feature_index_2[692] = 10'd352;
assign feature_index_2[693] = 10'd0;
assign feature_index_2[694] = 10'd0;
assign feature_index_2[695] = 10'd408;
assign feature_index_2[696] = 10'd513;
assign feature_index_2[697] = 10'd436;
assign feature_index_2[698] = 10'd267;
assign feature_index_2[699] = 10'd542;
assign feature_index_2[700] = 10'd547;
assign feature_index_2[701] = 10'd206;
assign feature_index_2[702] = 10'd272;
assign feature_index_2[703] = 10'd602;
assign feature_index_2[704] = 10'd318;
assign feature_index_2[705] = 10'd159;
assign feature_index_2[706] = 10'd509;
assign feature_index_2[707] = 10'd353;
assign feature_index_2[708] = 10'd539;
assign feature_index_2[709] = 10'd402;
assign feature_index_2[710] = 10'd156;
assign feature_index_2[711] = 10'd490;
assign feature_index_2[712] = 10'd185;
assign feature_index_2[713] = 10'd319;
assign feature_index_2[714] = 10'd606;
assign feature_index_2[715] = 10'd232;
assign feature_index_2[716] = 10'd274;
assign feature_index_2[717] = 10'd344;
assign feature_index_2[718] = 10'd638;
assign feature_index_2[719] = 10'd683;
assign feature_index_2[720] = 10'd554;
assign feature_index_2[721] = 10'd212;
assign feature_index_2[722] = 10'd568;
assign feature_index_2[723] = 10'd297;
assign feature_index_2[724] = 10'd592;
assign feature_index_2[725] = 10'd567;
assign feature_index_2[726] = 10'd0;
assign feature_index_2[727] = 10'd158;
assign feature_index_2[728] = 10'd295;
assign feature_index_2[729] = 10'd317;
assign feature_index_2[730] = 10'd470;
assign feature_index_2[731] = 10'd489;
assign feature_index_2[732] = 10'd467;
assign feature_index_2[733] = 10'd411;
assign feature_index_2[734] = 10'd575;
assign feature_index_2[735] = 10'd351;
assign feature_index_2[736] = 10'd0;
assign feature_index_2[737] = 10'd401;
assign feature_index_2[738] = 10'd0;
assign feature_index_2[739] = 10'd299;
assign feature_index_2[740] = 10'd522;
assign feature_index_2[741] = 10'd0;
assign feature_index_2[742] = 10'd0;
assign feature_index_2[743] = 10'd0;
assign feature_index_2[744] = 10'd0;
assign feature_index_2[745] = 10'd0;
assign feature_index_2[746] = 10'd0;
assign feature_index_2[747] = 10'd554;
assign feature_index_2[748] = 10'd101;
assign feature_index_2[749] = 10'd0;
assign feature_index_2[750] = 10'd0;
assign feature_index_2[751] = 10'd0;
assign feature_index_2[752] = 10'd0;
assign feature_index_2[753] = 10'd0;
assign feature_index_2[754] = 10'd0;
assign feature_index_2[755] = 10'd0;
assign feature_index_2[756] = 10'd0;
assign feature_index_2[757] = 10'd0;
assign feature_index_2[758] = 10'd0;
assign feature_index_2[759] = 10'd0;
assign feature_index_2[760] = 10'd0;
assign feature_index_2[761] = 10'd0;
assign feature_index_2[762] = 10'd0;
assign feature_index_2[763] = 10'd0;
assign feature_index_2[764] = 10'd0;
assign feature_index_2[765] = 10'd0;
assign feature_index_2[766] = 10'd0;
assign feature_index_2[767] = 10'd459;
assign feature_index_2[768] = 10'd236;
assign feature_index_2[769] = 10'd374;
assign feature_index_2[770] = 10'd0;
assign feature_index_2[771] = 10'd218;
assign feature_index_2[772] = 10'd354;
assign feature_index_2[773] = 10'd464;
assign feature_index_2[774] = 10'd373;
assign feature_index_2[775] = 10'd546;
assign feature_index_2[776] = 10'd0;
assign feature_index_2[777] = 10'd457;
assign feature_index_2[778] = 10'd0;
assign feature_index_2[779] = 10'd270;
assign feature_index_2[780] = 10'd221;
assign feature_index_2[781] = 10'd463;
assign feature_index_2[782] = 10'd267;
assign feature_index_2[783] = 10'd348;
assign feature_index_2[784] = 10'd174;
assign feature_index_2[785] = 10'd464;
assign feature_index_2[786] = 10'd0;
assign feature_index_2[787] = 10'd0;
assign feature_index_2[788] = 10'd0;
assign feature_index_2[789] = 10'd0;
assign feature_index_2[790] = 10'd0;
assign feature_index_2[791] = 10'd0;
assign feature_index_2[792] = 10'd0;
assign feature_index_2[793] = 10'd415;
assign feature_index_2[794] = 10'd275;
assign feature_index_2[795] = 10'd0;
assign feature_index_2[796] = 10'd0;
assign feature_index_2[797] = 10'd0;
assign feature_index_2[798] = 10'd0;
assign feature_index_2[799] = 10'd428;
assign feature_index_2[800] = 10'd680;
assign feature_index_2[801] = 10'd0;
assign feature_index_2[802] = 10'd204;
assign feature_index_2[803] = 10'd0;
assign feature_index_2[804] = 10'd180;
assign feature_index_2[805] = 10'd489;
assign feature_index_2[806] = 10'd456;
assign feature_index_2[807] = 10'd689;
assign feature_index_2[808] = 10'd0;
assign feature_index_2[809] = 10'd0;
assign feature_index_2[810] = 10'd0;
assign feature_index_2[811] = 10'd0;
assign feature_index_2[812] = 10'd594;
assign feature_index_2[813] = 10'd347;
assign feature_index_2[814] = 10'd0;
assign feature_index_2[815] = 10'd507;
assign feature_index_2[816] = 10'd0;
assign feature_index_2[817] = 10'd375;
assign feature_index_2[818] = 10'd0;
assign feature_index_2[819] = 10'd455;
assign feature_index_2[820] = 10'd425;
assign feature_index_2[821] = 10'd0;
assign feature_index_2[822] = 10'd130;
assign feature_index_2[823] = 10'd0;
assign feature_index_2[824] = 10'd540;
assign feature_index_2[825] = 10'd0;
assign feature_index_2[826] = 10'd375;
assign feature_index_2[827] = 10'd0;
assign feature_index_2[828] = 10'd239;
assign feature_index_2[829] = 10'd600;
assign feature_index_2[830] = 10'd156;
assign feature_index_2[831] = 10'd385;
assign feature_index_2[832] = 10'd411;
assign feature_index_2[833] = 10'd518;
assign feature_index_2[834] = 10'd0;
assign feature_index_2[835] = 10'd118;
assign feature_index_2[836] = 10'd682;
assign feature_index_2[837] = 10'd404;
assign feature_index_2[838] = 10'd0;
assign feature_index_2[839] = 10'd345;
assign feature_index_2[840] = 10'd664;
assign feature_index_2[841] = 10'd273;
assign feature_index_2[842] = 10'd215;
assign feature_index_2[843] = 10'd550;
assign feature_index_2[844] = 10'd594;
assign feature_index_2[845] = 10'd297;
assign feature_index_2[846] = 10'd659;
assign feature_index_2[847] = 10'd682;
assign feature_index_2[848] = 10'd520;
assign feature_index_2[849] = 10'd0;
assign feature_index_2[850] = 10'd515;
assign feature_index_2[851] = 10'd131;
assign feature_index_2[852] = 10'd0;
assign feature_index_2[853] = 10'd484;
assign feature_index_2[854] = 10'd547;
assign feature_index_2[855] = 10'd519;
assign feature_index_2[856] = 10'd405;
assign feature_index_2[857] = 10'd136;
assign feature_index_2[858] = 10'd243;
assign feature_index_2[859] = 10'd401;
assign feature_index_2[860] = 10'd291;
assign feature_index_2[861] = 10'd406;
assign feature_index_2[862] = 10'd0;
assign feature_index_2[863] = 10'd158;
assign feature_index_2[864] = 10'd189;
assign feature_index_2[865] = 10'd541;
assign feature_index_2[866] = 10'd432;
assign feature_index_2[867] = 10'd315;
assign feature_index_2[868] = 10'd296;
assign feature_index_2[869] = 10'd0;
assign feature_index_2[870] = 10'd0;
assign feature_index_2[871] = 10'd518;
assign feature_index_2[872] = 10'd332;
assign feature_index_2[873] = 10'd0;
assign feature_index_2[874] = 10'd0;
assign feature_index_2[875] = 10'd0;
assign feature_index_2[876] = 10'd0;
assign feature_index_2[877] = 10'd0;
assign feature_index_2[878] = 10'd0;
assign feature_index_2[879] = 10'd549;
assign feature_index_2[880] = 10'd301;
assign feature_index_2[881] = 10'd156;
assign feature_index_2[882] = 10'd434;
assign feature_index_2[883] = 10'd541;
assign feature_index_2[884] = 10'd706;
assign feature_index_2[885] = 10'd354;
assign feature_index_2[886] = 10'd545;
assign feature_index_2[887] = 10'd384;
assign feature_index_2[888] = 10'd0;
assign feature_index_2[889] = 10'd0;
assign feature_index_2[890] = 10'd0;
assign feature_index_2[891] = 10'd218;
assign feature_index_2[892] = 10'd180;
assign feature_index_2[893] = 10'd623;
assign feature_index_2[894] = 10'd665;
assign feature_index_2[895] = 10'd247;
assign feature_index_2[896] = 10'd348;
assign feature_index_2[897] = 10'd242;
assign feature_index_2[898] = 10'd270;
assign feature_index_2[899] = 10'd326;
assign feature_index_2[900] = 10'd612;
assign feature_index_2[901] = 10'd320;
assign feature_index_2[902] = 10'd343;
assign feature_index_2[903] = 10'd579;
assign feature_index_2[904] = 10'd541;
assign feature_index_2[905] = 10'd327;
assign feature_index_2[906] = 10'd271;
assign feature_index_2[907] = 10'd709;
assign feature_index_2[908] = 10'd297;
assign feature_index_2[909] = 10'd327;
assign feature_index_2[910] = 10'd513;
assign feature_index_2[911] = 10'd263;
assign feature_index_2[912] = 10'd240;
assign feature_index_2[913] = 10'd331;
assign feature_index_2[914] = 10'd0;
assign feature_index_2[915] = 10'd294;
assign feature_index_2[916] = 10'd350;
assign feature_index_2[917] = 10'd498;
assign feature_index_2[918] = 10'd593;
assign feature_index_2[919] = 10'd665;
assign feature_index_2[920] = 10'd427;
assign feature_index_2[921] = 10'd0;
assign feature_index_2[922] = 10'd0;
assign feature_index_2[923] = 10'd489;
assign feature_index_2[924] = 10'd482;
assign feature_index_2[925] = 10'd257;
assign feature_index_2[926] = 10'd98;
assign feature_index_2[927] = 10'd602;
assign feature_index_2[928] = 10'd181;
assign feature_index_2[929] = 10'd377;
assign feature_index_2[930] = 10'd0;
assign feature_index_2[931] = 10'd594;
assign feature_index_2[932] = 10'd707;
assign feature_index_2[933] = 10'd479;
assign feature_index_2[934] = 10'd234;
assign feature_index_2[935] = 10'd274;
assign feature_index_2[936] = 10'd95;
assign feature_index_2[937] = 10'd0;
assign feature_index_2[938] = 10'd404;
assign feature_index_2[939] = 10'd520;
assign feature_index_2[940] = 10'd347;
assign feature_index_2[941] = 10'd581;
assign feature_index_2[942] = 10'd357;
assign feature_index_2[943] = 10'd274;
assign feature_index_2[944] = 10'd0;
assign feature_index_2[945] = 10'd434;
assign feature_index_2[946] = 10'd0;
assign feature_index_2[947] = 10'd0;
assign feature_index_2[948] = 10'd467;
assign feature_index_2[949] = 10'd0;
assign feature_index_2[950] = 10'd0;
assign feature_index_2[951] = 10'd0;
assign feature_index_2[952] = 10'd378;
assign feature_index_2[953] = 10'd0;
assign feature_index_2[954] = 10'd356;
assign feature_index_2[955] = 10'd409;
assign feature_index_2[956] = 10'd403;
assign feature_index_2[957] = 10'd379;
assign feature_index_2[958] = 10'd598;
assign feature_index_2[959] = 10'd427;
assign feature_index_2[960] = 10'd160;
assign feature_index_2[961] = 10'd275;
assign feature_index_2[962] = 10'd373;
assign feature_index_2[963] = 10'd455;
assign feature_index_2[964] = 10'd270;
assign feature_index_2[965] = 10'd521;
assign feature_index_2[966] = 10'd270;
assign feature_index_2[967] = 10'd150;
assign feature_index_2[968] = 10'd273;
assign feature_index_2[969] = 10'd0;
assign feature_index_2[970] = 10'd0;
assign feature_index_2[971] = 10'd470;
assign feature_index_2[972] = 10'd0;
assign feature_index_2[973] = 10'd0;
assign feature_index_2[974] = 10'd0;
assign feature_index_2[975] = 10'd658;
assign feature_index_2[976] = 10'd599;
assign feature_index_2[977] = 10'd0;
assign feature_index_2[978] = 10'd496;
assign feature_index_2[979] = 10'd322;
assign feature_index_2[980] = 10'd269;
assign feature_index_2[981] = 10'd608;
assign feature_index_2[982] = 10'd294;
assign feature_index_2[983] = 10'd321;
assign feature_index_2[984] = 10'd577;
assign feature_index_2[985] = 10'd351;
assign feature_index_2[986] = 10'd572;
assign feature_index_2[987] = 10'd0;
assign feature_index_2[988] = 10'd0;
assign feature_index_2[989] = 10'd429;
assign feature_index_2[990] = 10'd458;
assign feature_index_2[991] = 10'd466;
assign feature_index_2[992] = 10'd631;
assign feature_index_2[993] = 10'd185;
assign feature_index_2[994] = 10'd606;
assign feature_index_2[995] = 10'd567;
assign feature_index_2[996] = 10'd433;
assign feature_index_2[997] = 10'd510;
assign feature_index_2[998] = 10'd268;
assign feature_index_2[999] = 10'd658;
assign feature_index_2[1000] = 10'd331;
assign feature_index_2[1001] = 10'd0;
assign feature_index_2[1002] = 10'd0;
assign feature_index_2[1003] = 10'd705;
assign feature_index_2[1004] = 10'd607;
assign feature_index_2[1005] = 10'd495;
assign feature_index_2[1006] = 10'd500;
assign feature_index_2[1007] = 10'd355;
assign feature_index_2[1008] = 10'd0;
assign feature_index_2[1009] = 10'd470;
assign feature_index_2[1010] = 10'd288;
assign feature_index_2[1011] = 10'd304;
assign feature_index_2[1012] = 10'd0;
assign feature_index_2[1013] = 10'd327;
assign feature_index_2[1014] = 10'd0;
assign feature_index_2[1015] = 10'd495;
assign feature_index_2[1016] = 10'd269;
assign feature_index_2[1017] = 10'd509;
assign feature_index_2[1018] = 10'd455;
assign feature_index_2[1019] = 10'd652;
assign feature_index_2[1020] = 10'd550;
assign feature_index_2[1021] = 10'd0;
assign feature_index_2[1022] = 10'd264;
assign feature_index_3[0] = 10'd154;
assign feature_index_3[1] = 10'd740;
assign feature_index_3[2] = 10'd377;
assign feature_index_3[3] = 10'd434;
assign feature_index_3[4] = 10'd401;
assign feature_index_3[5] = 10'd357;
assign feature_index_3[6] = 10'd375;
assign feature_index_3[7] = 10'd594;
assign feature_index_3[8] = 10'd464;
assign feature_index_3[9] = 10'd347;
assign feature_index_3[10] = 10'd217;
assign feature_index_3[11] = 10'd123;
assign feature_index_3[12] = 10'd489;
assign feature_index_3[13] = 10'd486;
assign feature_index_3[14] = 10'd460;
assign feature_index_3[15] = 10'd432;
assign feature_index_3[16] = 10'd412;
assign feature_index_3[17] = 10'd402;
assign feature_index_3[18] = 10'd539;
assign feature_index_3[19] = 10'd210;
assign feature_index_3[20] = 10'd289;
assign feature_index_3[21] = 10'd461;
assign feature_index_3[22] = 10'd347;
assign feature_index_3[23] = 10'd542;
assign feature_index_3[24] = 10'd460;
assign feature_index_3[25] = 10'd461;
assign feature_index_3[26] = 10'd442;
assign feature_index_3[27] = 10'd550;
assign feature_index_3[28] = 10'd656;
assign feature_index_3[29] = 10'd289;
assign feature_index_3[30] = 10'd289;
assign feature_index_3[31] = 10'd511;
assign feature_index_3[32] = 10'd571;
assign feature_index_3[33] = 10'd497;
assign feature_index_3[34] = 10'd291;
assign feature_index_3[35] = 10'd263;
assign feature_index_3[36] = 10'd514;
assign feature_index_3[37] = 10'd402;
assign feature_index_3[38] = 10'd460;
assign feature_index_3[39] = 10'd457;
assign feature_index_3[40] = 10'd344;
assign feature_index_3[41] = 10'd406;
assign feature_index_3[42] = 10'd294;
assign feature_index_3[43] = 10'd240;
assign feature_index_3[44] = 10'd232;
assign feature_index_3[45] = 10'd382;
assign feature_index_3[46] = 10'd460;
assign feature_index_3[47] = 10'd460;
assign feature_index_3[48] = 10'd185;
assign feature_index_3[49] = 10'd320;
assign feature_index_3[50] = 10'd596;
assign feature_index_3[51] = 10'd210;
assign feature_index_3[52] = 10'd463;
assign feature_index_3[53] = 10'd537;
assign feature_index_3[54] = 10'd187;
assign feature_index_3[55] = 10'd214;
assign feature_index_3[56] = 10'd262;
assign feature_index_3[57] = 10'd399;
assign feature_index_3[58] = 10'd173;
assign feature_index_3[59] = 10'd291;
assign feature_index_3[60] = 10'd301;
assign feature_index_3[61] = 10'd515;
assign feature_index_3[62] = 10'd429;
assign feature_index_3[63] = 10'd401;
assign feature_index_3[64] = 10'd386;
assign feature_index_3[65] = 10'd210;
assign feature_index_3[66] = 10'd486;
assign feature_index_3[67] = 10'd149;
assign feature_index_3[68] = 10'd627;
assign feature_index_3[69] = 10'd580;
assign feature_index_3[70] = 10'd345;
assign feature_index_3[71] = 10'd296;
assign feature_index_3[72] = 10'd656;
assign feature_index_3[73] = 10'd596;
assign feature_index_3[74] = 10'd629;
assign feature_index_3[75] = 10'd484;
assign feature_index_3[76] = 10'd183;
assign feature_index_3[77] = 10'd218;
assign feature_index_3[78] = 10'd439;
assign feature_index_3[79] = 10'd0;
assign feature_index_3[80] = 10'd318;
assign feature_index_3[81] = 10'd455;
assign feature_index_3[82] = 10'd233;
assign feature_index_3[83] = 10'd491;
assign feature_index_3[84] = 10'd714;
assign feature_index_3[85] = 10'd243;
assign feature_index_3[86] = 10'd210;
assign feature_index_3[87] = 10'd484;
assign feature_index_3[88] = 10'd379;
assign feature_index_3[89] = 10'd572;
assign feature_index_3[90] = 10'd344;
assign feature_index_3[91] = 10'd262;
assign feature_index_3[92] = 10'd210;
assign feature_index_3[93] = 10'd433;
assign feature_index_3[94] = 10'd688;
assign feature_index_3[95] = 10'd427;
assign feature_index_3[96] = 10'd567;
assign feature_index_3[97] = 10'd267;
assign feature_index_3[98] = 10'd567;
assign feature_index_3[99] = 10'd70;
assign feature_index_3[100] = 10'd402;
assign feature_index_3[101] = 10'd293;
assign feature_index_3[102] = 10'd346;
assign feature_index_3[103] = 10'd158;
assign feature_index_3[104] = 10'd435;
assign feature_index_3[105] = 10'd217;
assign feature_index_3[106] = 10'd319;
assign feature_index_3[107] = 10'd374;
assign feature_index_3[108] = 10'd332;
assign feature_index_3[109] = 10'd660;
assign feature_index_3[110] = 10'd316;
assign feature_index_3[111] = 10'd381;
assign feature_index_3[112] = 10'd521;
assign feature_index_3[113] = 10'd544;
assign feature_index_3[114] = 10'd488;
assign feature_index_3[115] = 10'd517;
assign feature_index_3[116] = 10'd271;
assign feature_index_3[117] = 10'd126;
assign feature_index_3[118] = 10'd490;
assign feature_index_3[119] = 10'd483;
assign feature_index_3[120] = 10'd457;
assign feature_index_3[121] = 10'd216;
assign feature_index_3[122] = 10'd331;
assign feature_index_3[123] = 10'd514;
assign feature_index_3[124] = 10'd214;
assign feature_index_3[125] = 10'd541;
assign feature_index_3[126] = 10'd413;
assign feature_index_3[127] = 10'd513;
assign feature_index_3[128] = 10'd299;
assign feature_index_3[129] = 10'd463;
assign feature_index_3[130] = 10'd568;
assign feature_index_3[131] = 10'd513;
assign feature_index_3[132] = 10'd625;
assign feature_index_3[133] = 10'd344;
assign feature_index_3[134] = 10'd654;
assign feature_index_3[135] = 10'd325;
assign feature_index_3[136] = 10'd568;
assign feature_index_3[137] = 10'd408;
assign feature_index_3[138] = 10'd443;
assign feature_index_3[139] = 10'd428;
assign feature_index_3[140] = 10'd380;
assign feature_index_3[141] = 10'd352;
assign feature_index_3[142] = 10'd379;
assign feature_index_3[143] = 10'd381;
assign feature_index_3[144] = 10'd371;
assign feature_index_3[145] = 10'd344;
assign feature_index_3[146] = 10'd523;
assign feature_index_3[147] = 10'd266;
assign feature_index_3[148] = 10'd247;
assign feature_index_3[149] = 10'd298;
assign feature_index_3[150] = 10'd605;
assign feature_index_3[151] = 10'd376;
assign feature_index_3[152] = 10'd470;
assign feature_index_3[153] = 10'd266;
assign feature_index_3[154] = 10'd382;
assign feature_index_3[155] = 10'd455;
assign feature_index_3[156] = 10'd326;
assign feature_index_3[157] = 10'd681;
assign feature_index_3[158] = 10'd212;
assign feature_index_3[159] = 10'd0;
assign feature_index_3[160] = 10'd0;
assign feature_index_3[161] = 10'd0;
assign feature_index_3[162] = 10'd0;
assign feature_index_3[163] = 10'd354;
assign feature_index_3[164] = 10'd232;
assign feature_index_3[165] = 10'd455;
assign feature_index_3[166] = 10'd371;
assign feature_index_3[167] = 10'd0;
assign feature_index_3[168] = 10'd262;
assign feature_index_3[169] = 10'd0;
assign feature_index_3[170] = 10'd490;
assign feature_index_3[171] = 10'd210;
assign feature_index_3[172] = 10'd491;
assign feature_index_3[173] = 10'd0;
assign feature_index_3[174] = 10'd460;
assign feature_index_3[175] = 10'd427;
assign feature_index_3[176] = 10'd0;
assign feature_index_3[177] = 10'd293;
assign feature_index_3[178] = 10'd232;
assign feature_index_3[179] = 10'd0;
assign feature_index_3[180] = 10'd241;
assign feature_index_3[181] = 10'd629;
assign feature_index_3[182] = 10'd328;
assign feature_index_3[183] = 10'd680;
assign feature_index_3[184] = 10'd212;
assign feature_index_3[185] = 10'd403;
assign feature_index_3[186] = 10'd206;
assign feature_index_3[187] = 10'd0;
assign feature_index_3[188] = 10'd430;
assign feature_index_3[189] = 10'd301;
assign feature_index_3[190] = 10'd0;
assign feature_index_3[191] = 10'd491;
assign feature_index_3[192] = 10'd626;
assign feature_index_3[193] = 10'd326;
assign feature_index_3[194] = 10'd354;
assign feature_index_3[195] = 10'd537;
assign feature_index_3[196] = 10'd401;
assign feature_index_3[197] = 10'd325;
assign feature_index_3[198] = 10'd463;
assign feature_index_3[199] = 10'd415;
assign feature_index_3[200] = 10'd0;
assign feature_index_3[201] = 10'd577;
assign feature_index_3[202] = 10'd415;
assign feature_index_3[203] = 10'd398;
assign feature_index_3[204] = 10'd632;
assign feature_index_3[205] = 10'd263;
assign feature_index_3[206] = 10'd546;
assign feature_index_3[207] = 10'd184;
assign feature_index_3[208] = 10'd349;
assign feature_index_3[209] = 10'd352;
assign feature_index_3[210] = 10'd158;
assign feature_index_3[211] = 10'd594;
assign feature_index_3[212] = 10'd0;
assign feature_index_3[213] = 10'd314;
assign feature_index_3[214] = 10'd512;
assign feature_index_3[215] = 10'd599;
assign feature_index_3[216] = 10'd216;
assign feature_index_3[217] = 10'd370;
assign feature_index_3[218] = 10'd441;
assign feature_index_3[219] = 10'd574;
assign feature_index_3[220] = 10'd540;
assign feature_index_3[221] = 10'd661;
assign feature_index_3[222] = 10'd300;
assign feature_index_3[223] = 10'd238;
assign feature_index_3[224] = 10'd267;
assign feature_index_3[225] = 10'd294;
assign feature_index_3[226] = 10'd263;
assign feature_index_3[227] = 10'd177;
assign feature_index_3[228] = 10'd547;
assign feature_index_3[229] = 10'd427;
assign feature_index_3[230] = 10'd659;
assign feature_index_3[231] = 10'd291;
assign feature_index_3[232] = 10'd373;
assign feature_index_3[233] = 10'd295;
assign feature_index_3[234] = 10'd186;
assign feature_index_3[235] = 10'd542;
assign feature_index_3[236] = 10'd151;
assign feature_index_3[237] = 10'd242;
assign feature_index_3[238] = 10'd0;
assign feature_index_3[239] = 10'd315;
assign feature_index_3[240] = 10'd631;
assign feature_index_3[241] = 10'd150;
assign feature_index_3[242] = 10'd379;
assign feature_index_3[243] = 10'd160;
assign feature_index_3[244] = 10'd270;
assign feature_index_3[245] = 10'd548;
assign feature_index_3[246] = 10'd208;
assign feature_index_3[247] = 10'd350;
assign feature_index_3[248] = 10'd264;
assign feature_index_3[249] = 10'd659;
assign feature_index_3[250] = 10'd125;
assign feature_index_3[251] = 10'd679;
assign feature_index_3[252] = 10'd346;
assign feature_index_3[253] = 10'd327;
assign feature_index_3[254] = 10'd270;
assign feature_index_3[255] = 10'd404;
assign feature_index_3[256] = 10'd398;
assign feature_index_3[257] = 10'd570;
assign feature_index_3[258] = 10'd486;
assign feature_index_3[259] = 10'd351;
assign feature_index_3[260] = 10'd597;
assign feature_index_3[261] = 10'd515;
assign feature_index_3[262] = 10'd243;
assign feature_index_3[263] = 10'd626;
assign feature_index_3[264] = 10'd316;
assign feature_index_3[265] = 10'd220;
assign feature_index_3[266] = 10'd485;
assign feature_index_3[267] = 10'd469;
assign feature_index_3[268] = 10'd539;
assign feature_index_3[269] = 10'd204;
assign feature_index_3[270] = 10'd257;
assign feature_index_3[271] = 10'd555;
assign feature_index_3[272] = 10'd185;
assign feature_index_3[273] = 10'd0;
assign feature_index_3[274] = 10'd0;
assign feature_index_3[275] = 10'd380;
assign feature_index_3[276] = 10'd210;
assign feature_index_3[277] = 10'd299;
assign feature_index_3[278] = 10'd302;
assign feature_index_3[279] = 10'd540;
assign feature_index_3[280] = 10'd294;
assign feature_index_3[281] = 10'd487;
assign feature_index_3[282] = 10'd257;
assign feature_index_3[283] = 10'd402;
assign feature_index_3[284] = 10'd183;
assign feature_index_3[285] = 10'd385;
assign feature_index_3[286] = 10'd510;
assign feature_index_3[287] = 10'd540;
assign feature_index_3[288] = 10'd293;
assign feature_index_3[289] = 10'd206;
assign feature_index_3[290] = 10'd148;
assign feature_index_3[291] = 10'd353;
assign feature_index_3[292] = 10'd414;
assign feature_index_3[293] = 10'd711;
assign feature_index_3[294] = 10'd353;
assign feature_index_3[295] = 10'd263;
assign feature_index_3[296] = 10'd148;
assign feature_index_3[297] = 10'd483;
assign feature_index_3[298] = 10'd356;
assign feature_index_3[299] = 10'd547;
assign feature_index_3[300] = 10'd523;
assign feature_index_3[301] = 10'd130;
assign feature_index_3[302] = 10'd495;
assign feature_index_3[303] = 10'd156;
assign feature_index_3[304] = 10'd570;
assign feature_index_3[305] = 10'd371;
assign feature_index_3[306] = 10'd371;
assign feature_index_3[307] = 10'd742;
assign feature_index_3[308] = 10'd353;
assign feature_index_3[309] = 10'd623;
assign feature_index_3[310] = 10'd571;
assign feature_index_3[311] = 10'd275;
assign feature_index_3[312] = 10'd385;
assign feature_index_3[313] = 10'd176;
assign feature_index_3[314] = 10'd413;
assign feature_index_3[315] = 10'd382;
assign feature_index_3[316] = 10'd488;
assign feature_index_3[317] = 10'd289;
assign feature_index_3[318] = 10'd658;
assign feature_index_3[319] = 10'd0;
assign feature_index_3[320] = 10'd0;
assign feature_index_3[321] = 10'd0;
assign feature_index_3[322] = 10'd0;
assign feature_index_3[323] = 10'd0;
assign feature_index_3[324] = 10'd0;
assign feature_index_3[325] = 10'd0;
assign feature_index_3[326] = 10'd0;
assign feature_index_3[327] = 10'd292;
assign feature_index_3[328] = 10'd437;
assign feature_index_3[329] = 10'd0;
assign feature_index_3[330] = 10'd0;
assign feature_index_3[331] = 10'd739;
assign feature_index_3[332] = 10'd0;
assign feature_index_3[333] = 10'd0;
assign feature_index_3[334] = 10'd456;
assign feature_index_3[335] = 10'd0;
assign feature_index_3[336] = 10'd0;
assign feature_index_3[337] = 10'd0;
assign feature_index_3[338] = 10'd348;
assign feature_index_3[339] = 10'd0;
assign feature_index_3[340] = 10'd0;
assign feature_index_3[341] = 10'd0;
assign feature_index_3[342] = 10'd0;
assign feature_index_3[343] = 10'd0;
assign feature_index_3[344] = 10'd437;
assign feature_index_3[345] = 10'd0;
assign feature_index_3[346] = 10'd350;
assign feature_index_3[347] = 10'd0;
assign feature_index_3[348] = 10'd0;
assign feature_index_3[349] = 10'd288;
assign feature_index_3[350] = 10'd655;
assign feature_index_3[351] = 10'd213;
assign feature_index_3[352] = 10'd234;
assign feature_index_3[353] = 10'd0;
assign feature_index_3[354] = 10'd0;
assign feature_index_3[355] = 10'd323;
assign feature_index_3[356] = 10'd320;
assign feature_index_3[357] = 10'd403;
assign feature_index_3[358] = 10'd431;
assign feature_index_3[359] = 10'd0;
assign feature_index_3[360] = 10'd0;
assign feature_index_3[361] = 10'd0;
assign feature_index_3[362] = 10'd300;
assign feature_index_3[363] = 10'd0;
assign feature_index_3[364] = 10'd0;
assign feature_index_3[365] = 10'd0;
assign feature_index_3[366] = 10'd496;
assign feature_index_3[367] = 10'd0;
assign feature_index_3[368] = 10'd0;
assign feature_index_3[369] = 10'd0;
assign feature_index_3[370] = 10'd0;
assign feature_index_3[371] = 10'd0;
assign feature_index_3[372] = 10'd269;
assign feature_index_3[373] = 10'd405;
assign feature_index_3[374] = 10'd490;
assign feature_index_3[375] = 10'd0;
assign feature_index_3[376] = 10'd0;
assign feature_index_3[377] = 10'd600;
assign feature_index_3[378] = 10'd212;
assign feature_index_3[379] = 10'd208;
assign feature_index_3[380] = 10'd0;
assign feature_index_3[381] = 10'd0;
assign feature_index_3[382] = 10'd0;
assign feature_index_3[383] = 10'd263;
assign feature_index_3[384] = 10'd325;
assign feature_index_3[385] = 10'd602;
assign feature_index_3[386] = 10'd431;
assign feature_index_3[387] = 10'd627;
assign feature_index_3[388] = 10'd486;
assign feature_index_3[389] = 10'd100;
assign feature_index_3[390] = 10'd379;
assign feature_index_3[391] = 10'd178;
assign feature_index_3[392] = 10'd345;
assign feature_index_3[393] = 10'd129;
assign feature_index_3[394] = 10'd462;
assign feature_index_3[395] = 10'd100;
assign feature_index_3[396] = 10'd411;
assign feature_index_3[397] = 10'd455;
assign feature_index_3[398] = 10'd298;
assign feature_index_3[399] = 10'd462;
assign feature_index_3[400] = 10'd435;
assign feature_index_3[401] = 10'd0;
assign feature_index_3[402] = 10'd0;
assign feature_index_3[403] = 10'd564;
assign feature_index_3[404] = 10'd234;
assign feature_index_3[405] = 10'd656;
assign feature_index_3[406] = 10'd0;
assign feature_index_3[407] = 10'd98;
assign feature_index_3[408] = 10'd261;
assign feature_index_3[409] = 10'd121;
assign feature_index_3[410] = 10'd456;
assign feature_index_3[411] = 10'd552;
assign feature_index_3[412] = 10'd437;
assign feature_index_3[413] = 10'd350;
assign feature_index_3[414] = 10'd163;
assign feature_index_3[415] = 10'd241;
assign feature_index_3[416] = 10'd295;
assign feature_index_3[417] = 10'd132;
assign feature_index_3[418] = 10'd683;
assign feature_index_3[419] = 10'd72;
assign feature_index_3[420] = 10'd343;
assign feature_index_3[421] = 10'd184;
assign feature_index_3[422] = 10'd535;
assign feature_index_3[423] = 10'd272;
assign feature_index_3[424] = 10'd683;
assign feature_index_3[425] = 10'd0;
assign feature_index_3[426] = 10'd0;
assign feature_index_3[427] = 10'd639;
assign feature_index_3[428] = 10'd624;
assign feature_index_3[429] = 10'd0;
assign feature_index_3[430] = 10'd629;
assign feature_index_3[431] = 10'd316;
assign feature_index_3[432] = 10'd387;
assign feature_index_3[433] = 10'd632;
assign feature_index_3[434] = 10'd522;
assign feature_index_3[435] = 10'd347;
assign feature_index_3[436] = 10'd292;
assign feature_index_3[437] = 10'd0;
assign feature_index_3[438] = 10'd0;
assign feature_index_3[439] = 10'd665;
assign feature_index_3[440] = 10'd270;
assign feature_index_3[441] = 10'd128;
assign feature_index_3[442] = 10'd315;
assign feature_index_3[443] = 10'd0;
assign feature_index_3[444] = 10'd570;
assign feature_index_3[445] = 10'd244;
assign feature_index_3[446] = 10'd440;
assign feature_index_3[447] = 10'd518;
assign feature_index_3[448] = 10'd149;
assign feature_index_3[449] = 10'd489;
assign feature_index_3[450] = 10'd438;
assign feature_index_3[451] = 10'd321;
assign feature_index_3[452] = 10'd268;
assign feature_index_3[453] = 10'd384;
assign feature_index_3[454] = 10'd174;
assign feature_index_3[455] = 10'd296;
assign feature_index_3[456] = 10'd480;
assign feature_index_3[457] = 10'd177;
assign feature_index_3[458] = 10'd567;
assign feature_index_3[459] = 10'd243;
assign feature_index_3[460] = 10'd245;
assign feature_index_3[461] = 10'd456;
assign feature_index_3[462] = 10'd538;
assign feature_index_3[463] = 10'd383;
assign feature_index_3[464] = 10'd400;
assign feature_index_3[465] = 10'd347;
assign feature_index_3[466] = 10'd0;
assign feature_index_3[467] = 10'd246;
assign feature_index_3[468] = 10'd663;
assign feature_index_3[469] = 10'd301;
assign feature_index_3[470] = 10'd479;
assign feature_index_3[471] = 10'd568;
assign feature_index_3[472] = 10'd664;
assign feature_index_3[473] = 10'd153;
assign feature_index_3[474] = 10'd293;
assign feature_index_3[475] = 10'd0;
assign feature_index_3[476] = 10'd542;
assign feature_index_3[477] = 10'd0;
assign feature_index_3[478] = 10'd0;
assign feature_index_3[479] = 10'd486;
assign feature_index_3[480] = 10'd270;
assign feature_index_3[481] = 10'd351;
assign feature_index_3[482] = 10'd428;
assign feature_index_3[483] = 10'd133;
assign feature_index_3[484] = 10'd215;
assign feature_index_3[485] = 10'd567;
assign feature_index_3[486] = 10'd100;
assign feature_index_3[487] = 10'd270;
assign feature_index_3[488] = 10'd490;
assign feature_index_3[489] = 10'd489;
assign feature_index_3[490] = 10'd240;
assign feature_index_3[491] = 10'd484;
assign feature_index_3[492] = 10'd155;
assign feature_index_3[493] = 10'd0;
assign feature_index_3[494] = 10'd212;
assign feature_index_3[495] = 10'd319;
assign feature_index_3[496] = 10'd681;
assign feature_index_3[497] = 10'd657;
assign feature_index_3[498] = 10'd245;
assign feature_index_3[499] = 10'd268;
assign feature_index_3[500] = 10'd300;
assign feature_index_3[501] = 10'd484;
assign feature_index_3[502] = 10'd319;
assign feature_index_3[503] = 10'd593;
assign feature_index_3[504] = 10'd385;
assign feature_index_3[505] = 10'd440;
assign feature_index_3[506] = 10'd472;
assign feature_index_3[507] = 10'd543;
assign feature_index_3[508] = 10'd513;
assign feature_index_3[509] = 10'd99;
assign feature_index_3[510] = 10'd548;
assign feature_index_3[511] = 10'd259;
assign feature_index_3[512] = 10'd547;
assign feature_index_3[513] = 10'd378;
assign feature_index_3[514] = 10'd573;
assign feature_index_3[515] = 10'd297;
assign feature_index_3[516] = 10'd658;
assign feature_index_3[517] = 10'd640;
assign feature_index_3[518] = 10'd465;
assign feature_index_3[519] = 10'd543;
assign feature_index_3[520] = 10'd230;
assign feature_index_3[521] = 10'd185;
assign feature_index_3[522] = 10'd188;
assign feature_index_3[523] = 10'd436;
assign feature_index_3[524] = 10'd381;
assign feature_index_3[525] = 10'd189;
assign feature_index_3[526] = 10'd102;
assign feature_index_3[527] = 10'd68;
assign feature_index_3[528] = 10'd358;
assign feature_index_3[529] = 10'd516;
assign feature_index_3[530] = 10'd265;
assign feature_index_3[531] = 10'd217;
assign feature_index_3[532] = 10'd0;
assign feature_index_3[533] = 10'd380;
assign feature_index_3[534] = 10'd296;
assign feature_index_3[535] = 10'd102;
assign feature_index_3[536] = 10'd202;
assign feature_index_3[537] = 10'd405;
assign feature_index_3[538] = 10'd406;
assign feature_index_3[539] = 10'd247;
assign feature_index_3[540] = 10'd208;
assign feature_index_3[541] = 10'd488;
assign feature_index_3[542] = 10'd0;
assign feature_index_3[543] = 10'd512;
assign feature_index_3[544] = 10'd656;
assign feature_index_3[545] = 10'd73;
assign feature_index_3[546] = 10'd162;
assign feature_index_3[547] = 10'd0;
assign feature_index_3[548] = 10'd0;
assign feature_index_3[549] = 10'd0;
assign feature_index_3[550] = 10'd0;
assign feature_index_3[551] = 10'd129;
assign feature_index_3[552] = 10'd0;
assign feature_index_3[553] = 10'd285;
assign feature_index_3[554] = 10'd0;
assign feature_index_3[555] = 10'd439;
assign feature_index_3[556] = 10'd580;
assign feature_index_3[557] = 10'd570;
assign feature_index_3[558] = 10'd304;
assign feature_index_3[559] = 10'd542;
assign feature_index_3[560] = 10'd380;
assign feature_index_3[561] = 10'd208;
assign feature_index_3[562] = 10'd494;
assign feature_index_3[563] = 10'd102;
assign feature_index_3[564] = 10'd0;
assign feature_index_3[565] = 10'd522;
assign feature_index_3[566] = 10'd0;
assign feature_index_3[567] = 10'd464;
assign feature_index_3[568] = 10'd626;
assign feature_index_3[569] = 10'd608;
assign feature_index_3[570] = 10'd353;
assign feature_index_3[571] = 10'd456;
assign feature_index_3[572] = 10'd461;
assign feature_index_3[573] = 10'd376;
assign feature_index_3[574] = 10'd377;
assign feature_index_3[575] = 10'd458;
assign feature_index_3[576] = 10'd301;
assign feature_index_3[577] = 10'd242;
assign feature_index_3[578] = 10'd522;
assign feature_index_3[579] = 10'd578;
assign feature_index_3[580] = 10'd551;
assign feature_index_3[581] = 10'd524;
assign feature_index_3[582] = 10'd0;
assign feature_index_3[583] = 10'd515;
assign feature_index_3[584] = 10'd552;
assign feature_index_3[585] = 10'd652;
assign feature_index_3[586] = 10'd610;
assign feature_index_3[587] = 10'd184;
assign feature_index_3[588] = 10'd328;
assign feature_index_3[589] = 10'd687;
assign feature_index_3[590] = 10'd347;
assign feature_index_3[591] = 10'd210;
assign feature_index_3[592] = 10'd97;
assign feature_index_3[593] = 10'd188;
assign feature_index_3[594] = 10'd316;
assign feature_index_3[595] = 10'd317;
assign feature_index_3[596] = 10'd495;
assign feature_index_3[597] = 10'd661;
assign feature_index_3[598] = 10'd379;
assign feature_index_3[599] = 10'd576;
assign feature_index_3[600] = 10'd625;
assign feature_index_3[601] = 10'd510;
assign feature_index_3[602] = 10'd599;
assign feature_index_3[603] = 10'd656;
assign feature_index_3[604] = 10'd133;
assign feature_index_3[605] = 10'd353;
assign feature_index_3[606] = 10'd172;
assign feature_index_3[607] = 10'd432;
assign feature_index_3[608] = 10'd517;
assign feature_index_3[609] = 10'd632;
assign feature_index_3[610] = 10'd576;
assign feature_index_3[611] = 10'd685;
assign feature_index_3[612] = 10'd149;
assign feature_index_3[613] = 10'd203;
assign feature_index_3[614] = 10'd570;
assign feature_index_3[615] = 10'd525;
assign feature_index_3[616] = 10'd216;
assign feature_index_3[617] = 10'd356;
assign feature_index_3[618] = 10'd267;
assign feature_index_3[619] = 10'd485;
assign feature_index_3[620] = 10'd324;
assign feature_index_3[621] = 10'd155;
assign feature_index_3[622] = 10'd576;
assign feature_index_3[623] = 10'd103;
assign feature_index_3[624] = 10'd0;
assign feature_index_3[625] = 10'd272;
assign feature_index_3[626] = 10'd640;
assign feature_index_3[627] = 10'd329;
assign feature_index_3[628] = 10'd376;
assign feature_index_3[629] = 10'd220;
assign feature_index_3[630] = 10'd0;
assign feature_index_3[631] = 10'd514;
assign feature_index_3[632] = 10'd481;
assign feature_index_3[633] = 10'd606;
assign feature_index_3[634] = 10'd408;
assign feature_index_3[635] = 10'd401;
assign feature_index_3[636] = 10'd598;
assign feature_index_3[637] = 10'd592;
assign feature_index_3[638] = 10'd360;
assign feature_index_3[639] = 10'd0;
assign feature_index_3[640] = 10'd0;
assign feature_index_3[641] = 10'd0;
assign feature_index_3[642] = 10'd0;
assign feature_index_3[643] = 10'd0;
assign feature_index_3[644] = 10'd0;
assign feature_index_3[645] = 10'd0;
assign feature_index_3[646] = 10'd0;
assign feature_index_3[647] = 10'd0;
assign feature_index_3[648] = 10'd0;
assign feature_index_3[649] = 10'd0;
assign feature_index_3[650] = 10'd0;
assign feature_index_3[651] = 10'd0;
assign feature_index_3[652] = 10'd0;
assign feature_index_3[653] = 10'd0;
assign feature_index_3[654] = 10'd0;
assign feature_index_3[655] = 10'd0;
assign feature_index_3[656] = 10'd263;
assign feature_index_3[657] = 10'd462;
assign feature_index_3[658] = 10'd378;
assign feature_index_3[659] = 10'd0;
assign feature_index_3[660] = 10'd0;
assign feature_index_3[661] = 10'd0;
assign feature_index_3[662] = 10'd0;
assign feature_index_3[663] = 10'd631;
assign feature_index_3[664] = 10'd0;
assign feature_index_3[665] = 10'd0;
assign feature_index_3[666] = 10'd0;
assign feature_index_3[667] = 10'd0;
assign feature_index_3[668] = 10'd0;
assign feature_index_3[669] = 10'd0;
assign feature_index_3[670] = 10'd0;
assign feature_index_3[671] = 10'd0;
assign feature_index_3[672] = 10'd0;
assign feature_index_3[673] = 10'd0;
assign feature_index_3[674] = 10'd0;
assign feature_index_3[675] = 10'd0;
assign feature_index_3[676] = 10'd0;
assign feature_index_3[677] = 10'd212;
assign feature_index_3[678] = 10'd346;
assign feature_index_3[679] = 10'd0;
assign feature_index_3[680] = 10'd0;
assign feature_index_3[681] = 10'd0;
assign feature_index_3[682] = 10'd0;
assign feature_index_3[683] = 10'd0;
assign feature_index_3[684] = 10'd0;
assign feature_index_3[685] = 10'd0;
assign feature_index_3[686] = 10'd0;
assign feature_index_3[687] = 10'd0;
assign feature_index_3[688] = 10'd0;
assign feature_index_3[689] = 10'd432;
assign feature_index_3[690] = 10'd0;
assign feature_index_3[691] = 10'd0;
assign feature_index_3[692] = 10'd0;
assign feature_index_3[693] = 10'd264;
assign feature_index_3[694] = 10'd0;
assign feature_index_3[695] = 10'd0;
assign feature_index_3[696] = 10'd0;
assign feature_index_3[697] = 10'd0;
assign feature_index_3[698] = 10'd0;
assign feature_index_3[699] = 10'd682;
assign feature_index_3[700] = 10'd466;
assign feature_index_3[701] = 10'd570;
assign feature_index_3[702] = 10'd0;
assign feature_index_3[703] = 10'd0;
assign feature_index_3[704] = 10'd382;
assign feature_index_3[705] = 10'd0;
assign feature_index_3[706] = 10'd577;
assign feature_index_3[707] = 10'd0;
assign feature_index_3[708] = 10'd0;
assign feature_index_3[709] = 10'd0;
assign feature_index_3[710] = 10'd0;
assign feature_index_3[711] = 10'd347;
assign feature_index_3[712] = 10'd686;
assign feature_index_3[713] = 10'd210;
assign feature_index_3[714] = 10'd0;
assign feature_index_3[715] = 10'd0;
assign feature_index_3[716] = 10'd457;
assign feature_index_3[717] = 10'd0;
assign feature_index_3[718] = 10'd203;
assign feature_index_3[719] = 10'd0;
assign feature_index_3[720] = 10'd0;
assign feature_index_3[721] = 10'd0;
assign feature_index_3[722] = 10'd0;
assign feature_index_3[723] = 10'd0;
assign feature_index_3[724] = 10'd0;
assign feature_index_3[725] = 10'd320;
assign feature_index_3[726] = 10'd459;
assign feature_index_3[727] = 10'd0;
assign feature_index_3[728] = 10'd0;
assign feature_index_3[729] = 10'd0;
assign feature_index_3[730] = 10'd0;
assign feature_index_3[731] = 10'd0;
assign feature_index_3[732] = 10'd0;
assign feature_index_3[733] = 10'd625;
assign feature_index_3[734] = 10'd0;
assign feature_index_3[735] = 10'd0;
assign feature_index_3[736] = 10'd0;
assign feature_index_3[737] = 10'd0;
assign feature_index_3[738] = 10'd0;
assign feature_index_3[739] = 10'd0;
assign feature_index_3[740] = 10'd0;
assign feature_index_3[741] = 10'd0;
assign feature_index_3[742] = 10'd0;
assign feature_index_3[743] = 10'd0;
assign feature_index_3[744] = 10'd0;
assign feature_index_3[745] = 10'd239;
assign feature_index_3[746] = 10'd0;
assign feature_index_3[747] = 10'd371;
assign feature_index_3[748] = 10'd0;
assign feature_index_3[749] = 10'd0;
assign feature_index_3[750] = 10'd273;
assign feature_index_3[751] = 10'd0;
assign feature_index_3[752] = 10'd0;
assign feature_index_3[753] = 10'd0;
assign feature_index_3[754] = 10'd0;
assign feature_index_3[755] = 10'd0;
assign feature_index_3[756] = 10'd0;
assign feature_index_3[757] = 10'd370;
assign feature_index_3[758] = 10'd0;
assign feature_index_3[759] = 10'd0;
assign feature_index_3[760] = 10'd0;
assign feature_index_3[761] = 10'd0;
assign feature_index_3[762] = 10'd0;
assign feature_index_3[763] = 10'd0;
assign feature_index_3[764] = 10'd0;
assign feature_index_3[765] = 10'd0;
assign feature_index_3[766] = 10'd0;
assign feature_index_3[767] = 10'd609;
assign feature_index_3[768] = 10'd325;
assign feature_index_3[769] = 10'd543;
assign feature_index_3[770] = 10'd270;
assign feature_index_3[771] = 10'd159;
assign feature_index_3[772] = 10'd0;
assign feature_index_3[773] = 10'd483;
assign feature_index_3[774] = 10'd482;
assign feature_index_3[775] = 10'd71;
assign feature_index_3[776] = 10'd269;
assign feature_index_3[777] = 10'd156;
assign feature_index_3[778] = 10'd288;
assign feature_index_3[779] = 10'd430;
assign feature_index_3[780] = 10'd0;
assign feature_index_3[781] = 10'd162;
assign feature_index_3[782] = 10'd684;
assign feature_index_3[783] = 10'd244;
assign feature_index_3[784] = 10'd400;
assign feature_index_3[785] = 10'd322;
assign feature_index_3[786] = 10'd245;
assign feature_index_3[787] = 10'd544;
assign feature_index_3[788] = 10'd298;
assign feature_index_3[789] = 10'd290;
assign feature_index_3[790] = 10'd271;
assign feature_index_3[791] = 10'd381;
assign feature_index_3[792] = 10'd209;
assign feature_index_3[793] = 10'd375;
assign feature_index_3[794] = 10'd467;
assign feature_index_3[795] = 10'd434;
assign feature_index_3[796] = 10'd351;
assign feature_index_3[797] = 10'd400;
assign feature_index_3[798] = 10'd302;
assign feature_index_3[799] = 10'd294;
assign feature_index_3[800] = 10'd342;
assign feature_index_3[801] = 10'd0;
assign feature_index_3[802] = 10'd0;
assign feature_index_3[803] = 10'd0;
assign feature_index_3[804] = 10'd0;
assign feature_index_3[805] = 10'd0;
assign feature_index_3[806] = 10'd0;
assign feature_index_3[807] = 10'd213;
assign feature_index_3[808] = 10'd0;
assign feature_index_3[809] = 10'd130;
assign feature_index_3[810] = 10'd487;
assign feature_index_3[811] = 10'd208;
assign feature_index_3[812] = 10'd428;
assign feature_index_3[813] = 10'd0;
assign feature_index_3[814] = 10'd0;
assign feature_index_3[815] = 10'd461;
assign feature_index_3[816] = 10'd70;
assign feature_index_3[817] = 10'd0;
assign feature_index_3[818] = 10'd471;
assign feature_index_3[819] = 10'd0;
assign feature_index_3[820] = 10'd0;
assign feature_index_3[821] = 10'd317;
assign feature_index_3[822] = 10'd409;
assign feature_index_3[823] = 10'd372;
assign feature_index_3[824] = 10'd0;
assign feature_index_3[825] = 10'd319;
assign feature_index_3[826] = 10'd570;
assign feature_index_3[827] = 10'd263;
assign feature_index_3[828] = 10'd0;
assign feature_index_3[829] = 10'd294;
assign feature_index_3[830] = 10'd0;
assign feature_index_3[831] = 10'd267;
assign feature_index_3[832] = 10'd320;
assign feature_index_3[833] = 10'd462;
assign feature_index_3[834] = 10'd455;
assign feature_index_3[835] = 10'd517;
assign feature_index_3[836] = 10'd571;
assign feature_index_3[837] = 10'd573;
assign feature_index_3[838] = 10'd0;
assign feature_index_3[839] = 10'd290;
assign feature_index_3[840] = 10'd0;
assign feature_index_3[841] = 10'd347;
assign feature_index_3[842] = 10'd174;
assign feature_index_3[843] = 10'd576;
assign feature_index_3[844] = 10'd242;
assign feature_index_3[845] = 10'd127;
assign feature_index_3[846] = 10'd0;
assign feature_index_3[847] = 10'd0;
assign feature_index_3[848] = 10'd0;
assign feature_index_3[849] = 10'd0;
assign feature_index_3[850] = 10'd0;
assign feature_index_3[851] = 10'd0;
assign feature_index_3[852] = 10'd0;
assign feature_index_3[853] = 10'd0;
assign feature_index_3[854] = 10'd0;
assign feature_index_3[855] = 10'd634;
assign feature_index_3[856] = 10'd287;
assign feature_index_3[857] = 10'd290;
assign feature_index_3[858] = 10'd0;
assign feature_index_3[859] = 10'd0;
assign feature_index_3[860] = 10'd0;
assign feature_index_3[861] = 10'd652;
assign feature_index_3[862] = 10'd0;
assign feature_index_3[863] = 10'd380;
assign feature_index_3[864] = 10'd213;
assign feature_index_3[865] = 10'd411;
assign feature_index_3[866] = 10'd483;
assign feature_index_3[867] = 10'd412;
assign feature_index_3[868] = 10'd206;
assign feature_index_3[869] = 10'd568;
assign feature_index_3[870] = 10'd179;
assign feature_index_3[871] = 10'd684;
assign feature_index_3[872] = 10'd635;
assign feature_index_3[873] = 10'd289;
assign feature_index_3[874] = 10'd0;
assign feature_index_3[875] = 10'd0;
assign feature_index_3[876] = 10'd0;
assign feature_index_3[877] = 10'd0;
assign feature_index_3[878] = 10'd0;
assign feature_index_3[879] = 10'd425;
assign feature_index_3[880] = 10'd499;
assign feature_index_3[881] = 10'd687;
assign feature_index_3[882] = 10'd214;
assign feature_index_3[883] = 10'd0;
assign feature_index_3[884] = 10'd0;
assign feature_index_3[885] = 10'd0;
assign feature_index_3[886] = 10'd629;
assign feature_index_3[887] = 10'd0;
assign feature_index_3[888] = 10'd0;
assign feature_index_3[889] = 10'd0;
assign feature_index_3[890] = 10'd0;
assign feature_index_3[891] = 10'd0;
assign feature_index_3[892] = 10'd455;
assign feature_index_3[893] = 10'd513;
assign feature_index_3[894] = 10'd423;
assign feature_index_3[895] = 10'd599;
assign feature_index_3[896] = 10'd599;
assign feature_index_3[897] = 10'd626;
assign feature_index_3[898] = 10'd172;
assign feature_index_3[899] = 10'd317;
assign feature_index_3[900] = 10'd126;
assign feature_index_3[901] = 10'd518;
assign feature_index_3[902] = 10'd607;
assign feature_index_3[903] = 10'd629;
assign feature_index_3[904] = 10'd651;
assign feature_index_3[905] = 10'd160;
assign feature_index_3[906] = 10'd595;
assign feature_index_3[907] = 10'd515;
assign feature_index_3[908] = 10'd0;
assign feature_index_3[909] = 10'd516;
assign feature_index_3[910] = 10'd0;
assign feature_index_3[911] = 10'd237;
assign feature_index_3[912] = 10'd155;
assign feature_index_3[913] = 10'd401;
assign feature_index_3[914] = 10'd178;
assign feature_index_3[915] = 10'd484;
assign feature_index_3[916] = 10'd461;
assign feature_index_3[917] = 10'd295;
assign feature_index_3[918] = 10'd489;
assign feature_index_3[919] = 10'd347;
assign feature_index_3[920] = 10'd319;
assign feature_index_3[921] = 10'd618;
assign feature_index_3[922] = 10'd358;
assign feature_index_3[923] = 10'd650;
assign feature_index_3[924] = 10'd0;
assign feature_index_3[925] = 10'd610;
assign feature_index_3[926] = 10'd322;
assign feature_index_3[927] = 10'd324;
assign feature_index_3[928] = 10'd403;
assign feature_index_3[929] = 10'd149;
assign feature_index_3[930] = 10'd213;
assign feature_index_3[931] = 10'd292;
assign feature_index_3[932] = 10'd261;
assign feature_index_3[933] = 10'd0;
assign feature_index_3[934] = 10'd0;
assign feature_index_3[935] = 10'd0;
assign feature_index_3[936] = 10'd0;
assign feature_index_3[937] = 10'd262;
assign feature_index_3[938] = 10'd385;
assign feature_index_3[939] = 10'd0;
assign feature_index_3[940] = 10'd184;
assign feature_index_3[941] = 10'd525;
assign feature_index_3[942] = 10'd0;
assign feature_index_3[943] = 10'd604;
assign feature_index_3[944] = 10'd523;
assign feature_index_3[945] = 10'd583;
assign feature_index_3[946] = 10'd610;
assign feature_index_3[947] = 10'd601;
assign feature_index_3[948] = 10'd129;
assign feature_index_3[949] = 10'd319;
assign feature_index_3[950] = 10'd554;
assign feature_index_3[951] = 10'd0;
assign feature_index_3[952] = 10'd0;
assign feature_index_3[953] = 10'd0;
assign feature_index_3[954] = 10'd0;
assign feature_index_3[955] = 10'd0;
assign feature_index_3[956] = 10'd0;
assign feature_index_3[957] = 10'd0;
assign feature_index_3[958] = 10'd0;
assign feature_index_3[959] = 10'd163;
assign feature_index_3[960] = 10'd459;
assign feature_index_3[961] = 10'd660;
assign feature_index_3[962] = 10'd412;
assign feature_index_3[963] = 10'd268;
assign feature_index_3[964] = 10'd628;
assign feature_index_3[965] = 10'd389;
assign feature_index_3[966] = 10'd121;
assign feature_index_3[967] = 10'd324;
assign feature_index_3[968] = 10'd212;
assign feature_index_3[969] = 10'd290;
assign feature_index_3[970] = 10'd388;
assign feature_index_3[971] = 10'd214;
assign feature_index_3[972] = 10'd101;
assign feature_index_3[973] = 10'd235;
assign feature_index_3[974] = 10'd538;
assign feature_index_3[975] = 10'd98;
assign feature_index_3[976] = 10'd650;
assign feature_index_3[977] = 10'd544;
assign feature_index_3[978] = 10'd206;
assign feature_index_3[979] = 10'd515;
assign feature_index_3[980] = 10'd316;
assign feature_index_3[981] = 10'd548;
assign feature_index_3[982] = 10'd517;
assign feature_index_3[983] = 10'd407;
assign feature_index_3[984] = 10'd174;
assign feature_index_3[985] = 10'd0;
assign feature_index_3[986] = 10'd265;
assign feature_index_3[987] = 10'd0;
assign feature_index_3[988] = 10'd0;
assign feature_index_3[989] = 10'd264;
assign feature_index_3[990] = 10'd272;
assign feature_index_3[991] = 10'd340;
assign feature_index_3[992] = 10'd299;
assign feature_index_3[993] = 10'd456;
assign feature_index_3[994] = 10'd539;
assign feature_index_3[995] = 10'd402;
assign feature_index_3[996] = 10'd371;
assign feature_index_3[997] = 10'd270;
assign feature_index_3[998] = 10'd459;
assign feature_index_3[999] = 10'd244;
assign feature_index_3[1000] = 10'd122;
assign feature_index_3[1001] = 10'd293;
assign feature_index_3[1002] = 10'd457;
assign feature_index_3[1003] = 10'd656;
assign feature_index_3[1004] = 10'd411;
assign feature_index_3[1005] = 10'd286;
assign feature_index_3[1006] = 10'd406;
assign feature_index_3[1007] = 10'd430;
assign feature_index_3[1008] = 10'd232;
assign feature_index_3[1009] = 10'd345;
assign feature_index_3[1010] = 10'd0;
assign feature_index_3[1011] = 10'd573;
assign feature_index_3[1012] = 10'd212;
assign feature_index_3[1013] = 10'd427;
assign feature_index_3[1014] = 10'd0;
assign feature_index_3[1015] = 10'd215;
assign feature_index_3[1016] = 10'd556;
assign feature_index_3[1017] = 10'd571;
assign feature_index_3[1018] = 10'd380;
assign feature_index_3[1019] = 10'd545;
assign feature_index_3[1020] = 10'd230;
assign feature_index_3[1021] = 10'd519;
assign feature_index_3[1022] = 10'd241;
assign feature_index_4[0] = 10'd155;
assign feature_index_4[1] = 10'd401;
assign feature_index_4[2] = 10'd545;
assign feature_index_4[3] = 10'd409;
assign feature_index_4[4] = 10'd275;
assign feature_index_4[5] = 10'd414;
assign feature_index_4[6] = 10'd242;
assign feature_index_4[7] = 10'd234;
assign feature_index_4[8] = 10'd540;
assign feature_index_4[9] = 10'd183;
assign feature_index_4[10] = 10'd330;
assign feature_index_4[11] = 10'd290;
assign feature_index_4[12] = 10'd274;
assign feature_index_4[13] = 10'd514;
assign feature_index_4[14] = 10'd373;
assign feature_index_4[15] = 10'd347;
assign feature_index_4[16] = 10'd470;
assign feature_index_4[17] = 10'd266;
assign feature_index_4[18] = 10'd653;
assign feature_index_4[19] = 10'd572;
assign feature_index_4[20] = 10'd189;
assign feature_index_4[21] = 10'd296;
assign feature_index_4[22] = 10'd538;
assign feature_index_4[23] = 10'd292;
assign feature_index_4[24] = 10'd351;
assign feature_index_4[25] = 10'd300;
assign feature_index_4[26] = 10'd404;
assign feature_index_4[27] = 10'd483;
assign feature_index_4[28] = 10'd318;
assign feature_index_4[29] = 10'd541;
assign feature_index_4[30] = 10'd435;
assign feature_index_4[31] = 10'd467;
assign feature_index_4[32] = 10'd380;
assign feature_index_4[33] = 10'd459;
assign feature_index_4[34] = 10'd425;
assign feature_index_4[35] = 10'd237;
assign feature_index_4[36] = 10'd261;
assign feature_index_4[37] = 10'd387;
assign feature_index_4[38] = 10'd487;
assign feature_index_4[39] = 10'd714;
assign feature_index_4[40] = 10'd577;
assign feature_index_4[41] = 10'd348;
assign feature_index_4[42] = 10'd302;
assign feature_index_4[43] = 10'd356;
assign feature_index_4[44] = 10'd735;
assign feature_index_4[45] = 10'd464;
assign feature_index_4[46] = 10'd320;
assign feature_index_4[47] = 10'd351;
assign feature_index_4[48] = 10'd180;
assign feature_index_4[49] = 10'd435;
assign feature_index_4[50] = 10'd273;
assign feature_index_4[51] = 10'd492;
assign feature_index_4[52] = 10'd484;
assign feature_index_4[53] = 10'd344;
assign feature_index_4[54] = 10'd496;
assign feature_index_4[55] = 10'd375;
assign feature_index_4[56] = 10'd291;
assign feature_index_4[57] = 10'd179;
assign feature_index_4[58] = 10'd684;
assign feature_index_4[59] = 10'd350;
assign feature_index_4[60] = 10'd321;
assign feature_index_4[61] = 10'd324;
assign feature_index_4[62] = 10'd126;
assign feature_index_4[63] = 10'd273;
assign feature_index_4[64] = 10'd486;
assign feature_index_4[65] = 10'd467;
assign feature_index_4[66] = 10'd433;
assign feature_index_4[67] = 10'd405;
assign feature_index_4[68] = 10'd376;
assign feature_index_4[69] = 10'd464;
assign feature_index_4[70] = 10'd405;
assign feature_index_4[71] = 10'd427;
assign feature_index_4[72] = 10'd432;
assign feature_index_4[73] = 10'd550;
assign feature_index_4[74] = 10'd375;
assign feature_index_4[75] = 10'd375;
assign feature_index_4[76] = 10'd430;
assign feature_index_4[77] = 10'd632;
assign feature_index_4[78] = 10'd324;
assign feature_index_4[79] = 10'd655;
assign feature_index_4[80] = 10'd187;
assign feature_index_4[81] = 10'd460;
assign feature_index_4[82] = 10'd217;
assign feature_index_4[83] = 10'd527;
assign feature_index_4[84] = 10'd570;
assign feature_index_4[85] = 10'd105;
assign feature_index_4[86] = 10'd380;
assign feature_index_4[87] = 10'd299;
assign feature_index_4[88] = 10'd242;
assign feature_index_4[89] = 10'd161;
assign feature_index_4[90] = 10'd208;
assign feature_index_4[91] = 10'd95;
assign feature_index_4[92] = 10'd242;
assign feature_index_4[93] = 10'd316;
assign feature_index_4[94] = 10'd461;
assign feature_index_4[95] = 10'd461;
assign feature_index_4[96] = 10'd515;
assign feature_index_4[97] = 10'd329;
assign feature_index_4[98] = 10'd179;
assign feature_index_4[99] = 10'd242;
assign feature_index_4[100] = 10'd102;
assign feature_index_4[101] = 10'd488;
assign feature_index_4[102] = 10'd541;
assign feature_index_4[103] = 10'd488;
assign feature_index_4[104] = 10'd568;
assign feature_index_4[105] = 10'd324;
assign feature_index_4[106] = 10'd437;
assign feature_index_4[107] = 10'd658;
assign feature_index_4[108] = 10'd600;
assign feature_index_4[109] = 10'd398;
assign feature_index_4[110] = 10'd291;
assign feature_index_4[111] = 10'd300;
assign feature_index_4[112] = 10'd262;
assign feature_index_4[113] = 10'd317;
assign feature_index_4[114] = 10'd625;
assign feature_index_4[115] = 10'd403;
assign feature_index_4[116] = 10'd400;
assign feature_index_4[117] = 10'd653;
assign feature_index_4[118] = 10'd399;
assign feature_index_4[119] = 10'd346;
assign feature_index_4[120] = 10'd651;
assign feature_index_4[121] = 10'd343;
assign feature_index_4[122] = 10'd609;
assign feature_index_4[123] = 10'd597;
assign feature_index_4[124] = 10'd379;
assign feature_index_4[125] = 10'd657;
assign feature_index_4[126] = 10'd455;
assign feature_index_4[127] = 10'd553;
assign feature_index_4[128] = 10'd377;
assign feature_index_4[129] = 10'd312;
assign feature_index_4[130] = 10'd607;
assign feature_index_4[131] = 10'd104;
assign feature_index_4[132] = 10'd341;
assign feature_index_4[133] = 10'd713;
assign feature_index_4[134] = 10'd161;
assign feature_index_4[135] = 10'd596;
assign feature_index_4[136] = 10'd488;
assign feature_index_4[137] = 10'd528;
assign feature_index_4[138] = 10'd528;
assign feature_index_4[139] = 10'd330;
assign feature_index_4[140] = 10'd600;
assign feature_index_4[141] = 10'd695;
assign feature_index_4[142] = 10'd461;
assign feature_index_4[143] = 10'd652;
assign feature_index_4[144] = 10'd207;
assign feature_index_4[145] = 10'd485;
assign feature_index_4[146] = 10'd315;
assign feature_index_4[147] = 10'd406;
assign feature_index_4[148] = 10'd487;
assign feature_index_4[149] = 10'd607;
assign feature_index_4[150] = 10'd546;
assign feature_index_4[151] = 10'd684;
assign feature_index_4[152] = 10'd459;
assign feature_index_4[153] = 10'd266;
assign feature_index_4[154] = 10'd574;
assign feature_index_4[155] = 10'd294;
assign feature_index_4[156] = 10'd185;
assign feature_index_4[157] = 10'd435;
assign feature_index_4[158] = 10'd245;
assign feature_index_4[159] = 10'd717;
assign feature_index_4[160] = 10'd382;
assign feature_index_4[161] = 10'd459;
assign feature_index_4[162] = 10'd266;
assign feature_index_4[163] = 10'd739;
assign feature_index_4[164] = 10'd540;
assign feature_index_4[165] = 10'd659;
assign feature_index_4[166] = 10'd491;
assign feature_index_4[167] = 10'd354;
assign feature_index_4[168] = 10'd489;
assign feature_index_4[169] = 10'd178;
assign feature_index_4[170] = 10'd326;
assign feature_index_4[171] = 10'd248;
assign feature_index_4[172] = 10'd602;
assign feature_index_4[173] = 10'd624;
assign feature_index_4[174] = 10'd516;
assign feature_index_4[175] = 10'd414;
assign feature_index_4[176] = 10'd519;
assign feature_index_4[177] = 10'd428;
assign feature_index_4[178] = 10'd437;
assign feature_index_4[179] = 10'd207;
assign feature_index_4[180] = 10'd432;
assign feature_index_4[181] = 10'd213;
assign feature_index_4[182] = 10'd0;
assign feature_index_4[183] = 10'd409;
assign feature_index_4[184] = 10'd0;
assign feature_index_4[185] = 10'd399;
assign feature_index_4[186] = 10'd633;
assign feature_index_4[187] = 10'd323;
assign feature_index_4[188] = 10'd461;
assign feature_index_4[189] = 10'd427;
assign feature_index_4[190] = 10'd382;
assign feature_index_4[191] = 10'd455;
assign feature_index_4[192] = 10'd568;
assign feature_index_4[193] = 10'd376;
assign feature_index_4[194] = 10'd317;
assign feature_index_4[195] = 10'd270;
assign feature_index_4[196] = 10'd432;
assign feature_index_4[197] = 10'd460;
assign feature_index_4[198] = 10'd149;
assign feature_index_4[199] = 10'd485;
assign feature_index_4[200] = 10'd462;
assign feature_index_4[201] = 10'd271;
assign feature_index_4[202] = 10'd182;
assign feature_index_4[203] = 10'd299;
assign feature_index_4[204] = 10'd655;
assign feature_index_4[205] = 10'd488;
assign feature_index_4[206] = 10'd433;
assign feature_index_4[207] = 10'd316;
assign feature_index_4[208] = 10'd297;
assign feature_index_4[209] = 10'd626;
assign feature_index_4[210] = 10'd385;
assign feature_index_4[211] = 10'd354;
assign feature_index_4[212] = 10'd651;
assign feature_index_4[213] = 10'd408;
assign feature_index_4[214] = 10'd522;
assign feature_index_4[215] = 10'd425;
assign feature_index_4[216] = 10'd379;
assign feature_index_4[217] = 10'd491;
assign feature_index_4[218] = 10'd0;
assign feature_index_4[219] = 10'd535;
assign feature_index_4[220] = 10'd550;
assign feature_index_4[221] = 10'd341;
assign feature_index_4[222] = 10'd353;
assign feature_index_4[223] = 10'd177;
assign feature_index_4[224] = 10'd407;
assign feature_index_4[225] = 10'd658;
assign feature_index_4[226] = 10'd567;
assign feature_index_4[227] = 10'd297;
assign feature_index_4[228] = 10'd161;
assign feature_index_4[229] = 10'd486;
assign feature_index_4[230] = 10'd100;
assign feature_index_4[231] = 10'd652;
assign feature_index_4[232] = 10'd300;
assign feature_index_4[233] = 10'd343;
assign feature_index_4[234] = 10'd217;
assign feature_index_4[235] = 10'd658;
assign feature_index_4[236] = 10'd433;
assign feature_index_4[237] = 10'd460;
assign feature_index_4[238] = 10'd297;
assign feature_index_4[239] = 10'd578;
assign feature_index_4[240] = 10'd293;
assign feature_index_4[241] = 10'd292;
assign feature_index_4[242] = 10'd248;
assign feature_index_4[243] = 10'd687;
assign feature_index_4[244] = 10'd492;
assign feature_index_4[245] = 10'd657;
assign feature_index_4[246] = 10'd514;
assign feature_index_4[247] = 10'd570;
assign feature_index_4[248] = 10'd211;
assign feature_index_4[249] = 10'd484;
assign feature_index_4[250] = 10'd515;
assign feature_index_4[251] = 10'd455;
assign feature_index_4[252] = 10'd441;
assign feature_index_4[253] = 10'd377;
assign feature_index_4[254] = 10'd481;
assign feature_index_4[255] = 10'd522;
assign feature_index_4[256] = 10'd300;
assign feature_index_4[257] = 10'd243;
assign feature_index_4[258] = 10'd248;
assign feature_index_4[259] = 10'd537;
assign feature_index_4[260] = 10'd0;
assign feature_index_4[261] = 10'd427;
assign feature_index_4[262] = 10'd349;
assign feature_index_4[263] = 10'd219;
assign feature_index_4[264] = 10'd570;
assign feature_index_4[265] = 10'd259;
assign feature_index_4[266] = 10'd554;
assign feature_index_4[267] = 10'd287;
assign feature_index_4[268] = 10'd548;
assign feature_index_4[269] = 10'd301;
assign feature_index_4[270] = 10'd510;
assign feature_index_4[271] = 10'd511;
assign feature_index_4[272] = 10'd399;
assign feature_index_4[273] = 10'd319;
assign feature_index_4[274] = 10'd348;
assign feature_index_4[275] = 10'd383;
assign feature_index_4[276] = 10'd0;
assign feature_index_4[277] = 10'd570;
assign feature_index_4[278] = 10'd125;
assign feature_index_4[279] = 10'd517;
assign feature_index_4[280] = 10'd379;
assign feature_index_4[281] = 10'd214;
assign feature_index_4[282] = 10'd240;
assign feature_index_4[283] = 10'd212;
assign feature_index_4[284] = 10'd0;
assign feature_index_4[285] = 10'd0;
assign feature_index_4[286] = 10'd265;
assign feature_index_4[287] = 10'd293;
assign feature_index_4[288] = 10'd205;
assign feature_index_4[289] = 10'd326;
assign feature_index_4[290] = 10'd241;
assign feature_index_4[291] = 10'd318;
assign feature_index_4[292] = 10'd246;
assign feature_index_4[293] = 10'd523;
assign feature_index_4[294] = 10'd319;
assign feature_index_4[295] = 10'd456;
assign feature_index_4[296] = 10'd292;
assign feature_index_4[297] = 10'd179;
assign feature_index_4[298] = 10'd297;
assign feature_index_4[299] = 10'd580;
assign feature_index_4[300] = 10'd455;
assign feature_index_4[301] = 10'd346;
assign feature_index_4[302] = 10'd551;
assign feature_index_4[303] = 10'd343;
assign feature_index_4[304] = 10'd634;
assign feature_index_4[305] = 10'd525;
assign feature_index_4[306] = 10'd157;
assign feature_index_4[307] = 10'd158;
assign feature_index_4[308] = 10'd525;
assign feature_index_4[309] = 10'd524;
assign feature_index_4[310] = 10'd318;
assign feature_index_4[311] = 10'd542;
assign feature_index_4[312] = 10'd312;
assign feature_index_4[313] = 10'd459;
assign feature_index_4[314] = 10'd347;
assign feature_index_4[315] = 10'd130;
assign feature_index_4[316] = 10'd376;
assign feature_index_4[317] = 10'd410;
assign feature_index_4[318] = 10'd211;
assign feature_index_4[319] = 10'd210;
assign feature_index_4[320] = 10'd237;
assign feature_index_4[321] = 10'd329;
assign feature_index_4[322] = 10'd464;
assign feature_index_4[323] = 10'd211;
assign feature_index_4[324] = 10'd205;
assign feature_index_4[325] = 10'd349;
assign feature_index_4[326] = 10'd432;
assign feature_index_4[327] = 10'd381;
assign feature_index_4[328] = 10'd406;
assign feature_index_4[329] = 10'd710;
assign feature_index_4[330] = 10'd325;
assign feature_index_4[331] = 10'd691;
assign feature_index_4[332] = 10'd489;
assign feature_index_4[333] = 10'd151;
assign feature_index_4[334] = 10'd107;
assign feature_index_4[335] = 10'd568;
assign feature_index_4[336] = 10'd480;
assign feature_index_4[337] = 10'd435;
assign feature_index_4[338] = 10'd655;
assign feature_index_4[339] = 10'd468;
assign feature_index_4[340] = 10'd158;
assign feature_index_4[341] = 10'd208;
assign feature_index_4[342] = 10'd204;
assign feature_index_4[343] = 10'd191;
assign feature_index_4[344] = 10'd300;
assign feature_index_4[345] = 10'd0;
assign feature_index_4[346] = 10'd239;
assign feature_index_4[347] = 10'd213;
assign feature_index_4[348] = 10'd240;
assign feature_index_4[349] = 10'd274;
assign feature_index_4[350] = 10'd632;
assign feature_index_4[351] = 10'd243;
assign feature_index_4[352] = 10'd0;
assign feature_index_4[353] = 10'd0;
assign feature_index_4[354] = 10'd606;
assign feature_index_4[355] = 10'd277;
assign feature_index_4[356] = 10'd269;
assign feature_index_4[357] = 10'd0;
assign feature_index_4[358] = 10'd631;
assign feature_index_4[359] = 10'd248;
assign feature_index_4[360] = 10'd487;
assign feature_index_4[361] = 10'd517;
assign feature_index_4[362] = 10'd157;
assign feature_index_4[363] = 10'd0;
assign feature_index_4[364] = 10'd219;
assign feature_index_4[365] = 10'd0;
assign feature_index_4[366] = 10'd0;
assign feature_index_4[367] = 10'd241;
assign feature_index_4[368] = 10'd439;
assign feature_index_4[369] = 10'd0;
assign feature_index_4[370] = 10'd0;
assign feature_index_4[371] = 10'd212;
assign feature_index_4[372] = 10'd322;
assign feature_index_4[373] = 10'd430;
assign feature_index_4[374] = 10'd207;
assign feature_index_4[375] = 10'd627;
assign feature_index_4[376] = 10'd357;
assign feature_index_4[377] = 10'd353;
assign feature_index_4[378] = 10'd184;
assign feature_index_4[379] = 10'd516;
assign feature_index_4[380] = 10'd124;
assign feature_index_4[381] = 10'd385;
assign feature_index_4[382] = 10'd627;
assign feature_index_4[383] = 10'd323;
assign feature_index_4[384] = 10'd405;
assign feature_index_4[385] = 10'd659;
assign feature_index_4[386] = 10'd316;
assign feature_index_4[387] = 10'd326;
assign feature_index_4[388] = 10'd261;
assign feature_index_4[389] = 10'd488;
assign feature_index_4[390] = 10'd341;
assign feature_index_4[391] = 10'd187;
assign feature_index_4[392] = 10'd346;
assign feature_index_4[393] = 10'd466;
assign feature_index_4[394] = 10'd491;
assign feature_index_4[395] = 10'd327;
assign feature_index_4[396] = 10'd406;
assign feature_index_4[397] = 10'd543;
assign feature_index_4[398] = 10'd500;
assign feature_index_4[399] = 10'd372;
assign feature_index_4[400] = 10'd384;
assign feature_index_4[401] = 10'd650;
assign feature_index_4[402] = 10'd596;
assign feature_index_4[403] = 10'd300;
assign feature_index_4[404] = 10'd571;
assign feature_index_4[405] = 10'd0;
assign feature_index_4[406] = 10'd625;
assign feature_index_4[407] = 10'd159;
assign feature_index_4[408] = 10'd550;
assign feature_index_4[409] = 10'd154;
assign feature_index_4[410] = 10'd601;
assign feature_index_4[411] = 10'd483;
assign feature_index_4[412] = 10'd430;
assign feature_index_4[413] = 10'd572;
assign feature_index_4[414] = 10'd510;
assign feature_index_4[415] = 10'd296;
assign feature_index_4[416] = 10'd458;
assign feature_index_4[417] = 10'd661;
assign feature_index_4[418] = 10'd373;
assign feature_index_4[419] = 10'd238;
assign feature_index_4[420] = 10'd681;
assign feature_index_4[421] = 10'd631;
assign feature_index_4[422] = 10'd187;
assign feature_index_4[423] = 10'd498;
assign feature_index_4[424] = 10'd601;
assign feature_index_4[425] = 10'd342;
assign feature_index_4[426] = 10'd355;
assign feature_index_4[427] = 10'd428;
assign feature_index_4[428] = 10'd376;
assign feature_index_4[429] = 10'd652;
assign feature_index_4[430] = 10'd344;
assign feature_index_4[431] = 10'd320;
assign feature_index_4[432] = 10'd0;
assign feature_index_4[433] = 10'd0;
assign feature_index_4[434] = 10'd517;
assign feature_index_4[435] = 10'd0;
assign feature_index_4[436] = 10'd187;
assign feature_index_4[437] = 10'd0;
assign feature_index_4[438] = 10'd0;
assign feature_index_4[439] = 10'd147;
assign feature_index_4[440] = 10'd0;
assign feature_index_4[441] = 10'd0;
assign feature_index_4[442] = 10'd627;
assign feature_index_4[443] = 10'd298;
assign feature_index_4[444] = 10'd683;
assign feature_index_4[445] = 10'd518;
assign feature_index_4[446] = 10'd682;
assign feature_index_4[447] = 10'd439;
assign feature_index_4[448] = 10'd543;
assign feature_index_4[449] = 10'd325;
assign feature_index_4[450] = 10'd621;
assign feature_index_4[451] = 10'd265;
assign feature_index_4[452] = 10'd467;
assign feature_index_4[453] = 10'd682;
assign feature_index_4[454] = 10'd245;
assign feature_index_4[455] = 10'd360;
assign feature_index_4[456] = 10'd124;
assign feature_index_4[457] = 10'd243;
assign feature_index_4[458] = 10'd521;
assign feature_index_4[459] = 10'd682;
assign feature_index_4[460] = 10'd129;
assign feature_index_4[461] = 10'd433;
assign feature_index_4[462] = 10'd408;
assign feature_index_4[463] = 10'd655;
assign feature_index_4[464] = 10'd522;
assign feature_index_4[465] = 10'd296;
assign feature_index_4[466] = 10'd492;
assign feature_index_4[467] = 10'd686;
assign feature_index_4[468] = 10'd635;
assign feature_index_4[469] = 10'd399;
assign feature_index_4[470] = 10'd371;
assign feature_index_4[471] = 10'd595;
assign feature_index_4[472] = 10'd571;
assign feature_index_4[473] = 10'd358;
assign feature_index_4[474] = 10'd294;
assign feature_index_4[475] = 10'd496;
assign feature_index_4[476] = 10'd413;
assign feature_index_4[477] = 10'd0;
assign feature_index_4[478] = 10'd413;
assign feature_index_4[479] = 10'd348;
assign feature_index_4[480] = 10'd690;
assign feature_index_4[481] = 10'd659;
assign feature_index_4[482] = 10'd662;
assign feature_index_4[483] = 10'd523;
assign feature_index_4[484] = 10'd687;
assign feature_index_4[485] = 10'd297;
assign feature_index_4[486] = 10'd486;
assign feature_index_4[487] = 10'd150;
assign feature_index_4[488] = 10'd635;
assign feature_index_4[489] = 10'd627;
assign feature_index_4[490] = 10'd399;
assign feature_index_4[491] = 10'd629;
assign feature_index_4[492] = 10'd489;
assign feature_index_4[493] = 10'd239;
assign feature_index_4[494] = 10'd486;
assign feature_index_4[495] = 10'd686;
assign feature_index_4[496] = 10'd485;
assign feature_index_4[497] = 10'd609;
assign feature_index_4[498] = 10'd278;
assign feature_index_4[499] = 10'd210;
assign feature_index_4[500] = 10'd329;
assign feature_index_4[501] = 10'd264;
assign feature_index_4[502] = 10'd528;
assign feature_index_4[503] = 10'd567;
assign feature_index_4[504] = 10'd104;
assign feature_index_4[505] = 10'd687;
assign feature_index_4[506] = 10'd551;
assign feature_index_4[507] = 10'd661;
assign feature_index_4[508] = 10'd624;
assign feature_index_4[509] = 10'd218;
assign feature_index_4[510] = 10'd172;
assign feature_index_4[511] = 10'd147;
assign feature_index_4[512] = 10'd294;
assign feature_index_4[513] = 10'd658;
assign feature_index_4[514] = 10'd483;
assign feature_index_4[515] = 10'd463;
assign feature_index_4[516] = 10'd453;
assign feature_index_4[517] = 10'd242;
assign feature_index_4[518] = 10'd428;
assign feature_index_4[519] = 10'd291;
assign feature_index_4[520] = 10'd349;
assign feature_index_4[521] = 10'd0;
assign feature_index_4[522] = 10'd0;
assign feature_index_4[523] = 10'd244;
assign feature_index_4[524] = 10'd555;
assign feature_index_4[525] = 10'd594;
assign feature_index_4[526] = 10'd0;
assign feature_index_4[527] = 10'd177;
assign feature_index_4[528] = 10'd443;
assign feature_index_4[529] = 10'd0;
assign feature_index_4[530] = 10'd0;
assign feature_index_4[531] = 10'd397;
assign feature_index_4[532] = 10'd527;
assign feature_index_4[533] = 10'd539;
assign feature_index_4[534] = 10'd0;
assign feature_index_4[535] = 10'd150;
assign feature_index_4[536] = 10'd173;
assign feature_index_4[537] = 10'd211;
assign feature_index_4[538] = 10'd288;
assign feature_index_4[539] = 10'd487;
assign feature_index_4[540] = 10'd265;
assign feature_index_4[541] = 10'd382;
assign feature_index_4[542] = 10'd511;
assign feature_index_4[543] = 10'd150;
assign feature_index_4[544] = 10'd237;
assign feature_index_4[545] = 10'd323;
assign feature_index_4[546] = 10'd410;
assign feature_index_4[547] = 10'd208;
assign feature_index_4[548] = 10'd215;
assign feature_index_4[549] = 10'd610;
assign feature_index_4[550] = 10'd686;
assign feature_index_4[551] = 10'd405;
assign feature_index_4[552] = 10'd275;
assign feature_index_4[553] = 10'd0;
assign feature_index_4[554] = 10'd0;
assign feature_index_4[555] = 10'd383;
assign feature_index_4[556] = 10'd122;
assign feature_index_4[557] = 10'd0;
assign feature_index_4[558] = 10'd439;
assign feature_index_4[559] = 10'd521;
assign feature_index_4[560] = 10'd124;
assign feature_index_4[561] = 10'd411;
assign feature_index_4[562] = 10'd240;
assign feature_index_4[563] = 10'd217;
assign feature_index_4[564] = 10'd210;
assign feature_index_4[565] = 10'd246;
assign feature_index_4[566] = 10'd96;
assign feature_index_4[567] = 10'd359;
assign feature_index_4[568] = 10'd668;
assign feature_index_4[569] = 10'd0;
assign feature_index_4[570] = 10'd0;
assign feature_index_4[571] = 10'd0;
assign feature_index_4[572] = 10'd0;
assign feature_index_4[573] = 10'd340;
assign feature_index_4[574] = 10'd488;
assign feature_index_4[575] = 10'd297;
assign feature_index_4[576] = 10'd382;
assign feature_index_4[577] = 10'd209;
assign feature_index_4[578] = 10'd235;
assign feature_index_4[579] = 10'd573;
assign feature_index_4[580] = 10'd488;
assign feature_index_4[581] = 10'd183;
assign feature_index_4[582] = 10'd188;
assign feature_index_4[583] = 10'd349;
assign feature_index_4[584] = 10'd378;
assign feature_index_4[585] = 10'd597;
assign feature_index_4[586] = 10'd181;
assign feature_index_4[587] = 10'd318;
assign feature_index_4[588] = 10'd292;
assign feature_index_4[589] = 10'd598;
assign feature_index_4[590] = 10'd456;
assign feature_index_4[591] = 10'd298;
assign feature_index_4[592] = 10'd511;
assign feature_index_4[593] = 10'd462;
assign feature_index_4[594] = 10'd376;
assign feature_index_4[595] = 10'd340;
assign feature_index_4[596] = 10'd466;
assign feature_index_4[597] = 10'd405;
assign feature_index_4[598] = 10'd319;
assign feature_index_4[599] = 10'd595;
assign feature_index_4[600] = 10'd600;
assign feature_index_4[601] = 10'd460;
assign feature_index_4[602] = 10'd444;
assign feature_index_4[603] = 10'd399;
assign feature_index_4[604] = 10'd183;
assign feature_index_4[605] = 10'd298;
assign feature_index_4[606] = 10'd406;
assign feature_index_4[607] = 10'd461;
assign feature_index_4[608] = 10'd525;
assign feature_index_4[609] = 10'd373;
assign feature_index_4[610] = 10'd265;
assign feature_index_4[611] = 10'd210;
assign feature_index_4[612] = 10'd120;
assign feature_index_4[613] = 10'd331;
assign feature_index_4[614] = 10'd357;
assign feature_index_4[615] = 10'd690;
assign feature_index_4[616] = 10'd152;
assign feature_index_4[617] = 10'd400;
assign feature_index_4[618] = 10'd327;
assign feature_index_4[619] = 10'd457;
assign feature_index_4[620] = 10'd0;
assign feature_index_4[621] = 10'd0;
assign feature_index_4[622] = 10'd0;
assign feature_index_4[623] = 10'd431;
assign feature_index_4[624] = 10'd0;
assign feature_index_4[625] = 10'd355;
assign feature_index_4[626] = 10'd0;
assign feature_index_4[627] = 10'd215;
assign feature_index_4[628] = 10'd0;
assign feature_index_4[629] = 10'd266;
assign feature_index_4[630] = 10'd174;
assign feature_index_4[631] = 10'd0;
assign feature_index_4[632] = 10'd0;
assign feature_index_4[633] = 10'd465;
assign feature_index_4[634] = 10'd0;
assign feature_index_4[635] = 10'd602;
assign feature_index_4[636] = 10'd187;
assign feature_index_4[637] = 10'd629;
assign feature_index_4[638] = 10'd575;
assign feature_index_4[639] = 10'd740;
assign feature_index_4[640] = 10'd240;
assign feature_index_4[641] = 10'd380;
assign feature_index_4[642] = 10'd202;
assign feature_index_4[643] = 10'd219;
assign feature_index_4[644] = 10'd495;
assign feature_index_4[645] = 10'd488;
assign feature_index_4[646] = 10'd210;
assign feature_index_4[647] = 10'd376;
assign feature_index_4[648] = 10'd402;
assign feature_index_4[649] = 10'd240;
assign feature_index_4[650] = 10'd246;
assign feature_index_4[651] = 10'd0;
assign feature_index_4[652] = 10'd713;
assign feature_index_4[653] = 10'd547;
assign feature_index_4[654] = 10'd325;
assign feature_index_4[655] = 10'd406;
assign feature_index_4[656] = 10'd266;
assign feature_index_4[657] = 10'd378;
assign feature_index_4[658] = 10'd316;
assign feature_index_4[659] = 10'd399;
assign feature_index_4[660] = 10'd495;
assign feature_index_4[661] = 10'd546;
assign feature_index_4[662] = 10'd568;
assign feature_index_4[663] = 10'd285;
assign feature_index_4[664] = 10'd176;
assign feature_index_4[665] = 10'd290;
assign feature_index_4[666] = 10'd467;
assign feature_index_4[667] = 10'd384;
assign feature_index_4[668] = 10'd434;
assign feature_index_4[669] = 10'd626;
assign feature_index_4[670] = 10'd0;
assign feature_index_4[671] = 10'd548;
assign feature_index_4[672] = 10'd435;
assign feature_index_4[673] = 10'd519;
assign feature_index_4[674] = 10'd0;
assign feature_index_4[675] = 10'd350;
assign feature_index_4[676] = 10'd483;
assign feature_index_4[677] = 10'd386;
assign feature_index_4[678] = 10'd466;
assign feature_index_4[679] = 10'd210;
assign feature_index_4[680] = 10'd458;
assign feature_index_4[681] = 10'd262;
assign feature_index_4[682] = 10'd516;
assign feature_index_4[683] = 10'd150;
assign feature_index_4[684] = 10'd289;
assign feature_index_4[685] = 10'd484;
assign feature_index_4[686] = 10'd314;
assign feature_index_4[687] = 10'd300;
assign feature_index_4[688] = 10'd353;
assign feature_index_4[689] = 10'd385;
assign feature_index_4[690] = 10'd489;
assign feature_index_4[691] = 10'd0;
assign feature_index_4[692] = 10'd0;
assign feature_index_4[693] = 10'd0;
assign feature_index_4[694] = 10'd301;
assign feature_index_4[695] = 10'd0;
assign feature_index_4[696] = 10'd349;
assign feature_index_4[697] = 10'd0;
assign feature_index_4[698] = 10'd177;
assign feature_index_4[699] = 10'd0;
assign feature_index_4[700] = 10'd343;
assign feature_index_4[701] = 10'd514;
assign feature_index_4[702] = 10'd495;
assign feature_index_4[703] = 10'd320;
assign feature_index_4[704] = 10'd353;
assign feature_index_4[705] = 10'd0;
assign feature_index_4[706] = 10'd0;
assign feature_index_4[707] = 10'd0;
assign feature_index_4[708] = 10'd0;
assign feature_index_4[709] = 10'd354;
assign feature_index_4[710] = 10'd0;
assign feature_index_4[711] = 10'd236;
assign feature_index_4[712] = 10'd0;
assign feature_index_4[713] = 10'd184;
assign feature_index_4[714] = 10'd0;
assign feature_index_4[715] = 10'd0;
assign feature_index_4[716] = 10'd0;
assign feature_index_4[717] = 10'd654;
assign feature_index_4[718] = 10'd439;
assign feature_index_4[719] = 10'd410;
assign feature_index_4[720] = 10'd313;
assign feature_index_4[721] = 10'd623;
assign feature_index_4[722] = 10'd352;
assign feature_index_4[723] = 10'd464;
assign feature_index_4[724] = 10'd655;
assign feature_index_4[725] = 10'd456;
assign feature_index_4[726] = 10'd0;
assign feature_index_4[727] = 10'd0;
assign feature_index_4[728] = 10'd0;
assign feature_index_4[729] = 10'd0;
assign feature_index_4[730] = 10'd459;
assign feature_index_4[731] = 10'd0;
assign feature_index_4[732] = 10'd0;
assign feature_index_4[733] = 10'd0;
assign feature_index_4[734] = 10'd0;
assign feature_index_4[735] = 10'd292;
assign feature_index_4[736] = 10'd352;
assign feature_index_4[737] = 10'd495;
assign feature_index_4[738] = 10'd600;
assign feature_index_4[739] = 10'd0;
assign feature_index_4[740] = 10'd0;
assign feature_index_4[741] = 10'd0;
assign feature_index_4[742] = 10'd0;
assign feature_index_4[743] = 10'd465;
assign feature_index_4[744] = 10'd293;
assign feature_index_4[745] = 10'd388;
assign feature_index_4[746] = 10'd323;
assign feature_index_4[747] = 10'd371;
assign feature_index_4[748] = 10'd487;
assign feature_index_4[749] = 10'd244;
assign feature_index_4[750] = 10'd581;
assign feature_index_4[751] = 10'd124;
assign feature_index_4[752] = 10'd549;
assign feature_index_4[753] = 10'd0;
assign feature_index_4[754] = 10'd0;
assign feature_index_4[755] = 10'd352;
assign feature_index_4[756] = 10'd631;
assign feature_index_4[757] = 10'd459;
assign feature_index_4[758] = 10'd0;
assign feature_index_4[759] = 10'd435;
assign feature_index_4[760] = 10'd324;
assign feature_index_4[761] = 10'd372;
assign feature_index_4[762] = 10'd209;
assign feature_index_4[763] = 10'd579;
assign feature_index_4[764] = 10'd164;
assign feature_index_4[765] = 10'd508;
assign feature_index_4[766] = 10'd468;
assign feature_index_4[767] = 10'd660;
assign feature_index_4[768] = 10'd572;
assign feature_index_4[769] = 10'd572;
assign feature_index_4[770] = 10'd470;
assign feature_index_4[771] = 10'd541;
assign feature_index_4[772] = 10'd323;
assign feature_index_4[773] = 10'd319;
assign feature_index_4[774] = 10'd403;
assign feature_index_4[775] = 10'd429;
assign feature_index_4[776] = 10'd344;
assign feature_index_4[777] = 10'd314;
assign feature_index_4[778] = 10'd514;
assign feature_index_4[779] = 10'd431;
assign feature_index_4[780] = 10'd228;
assign feature_index_4[781] = 10'd405;
assign feature_index_4[782] = 10'd665;
assign feature_index_4[783] = 10'd571;
assign feature_index_4[784] = 10'd402;
assign feature_index_4[785] = 10'd550;
assign feature_index_4[786] = 10'd461;
assign feature_index_4[787] = 10'd376;
assign feature_index_4[788] = 10'd0;
assign feature_index_4[789] = 10'd462;
assign feature_index_4[790] = 10'd187;
assign feature_index_4[791] = 10'd514;
assign feature_index_4[792] = 10'd357;
assign feature_index_4[793] = 10'd427;
assign feature_index_4[794] = 10'd467;
assign feature_index_4[795] = 10'd458;
assign feature_index_4[796] = 10'd434;
assign feature_index_4[797] = 10'd319;
assign feature_index_4[798] = 10'd0;
assign feature_index_4[799] = 10'd241;
assign feature_index_4[800] = 10'd661;
assign feature_index_4[801] = 10'd657;
assign feature_index_4[802] = 10'd349;
assign feature_index_4[803] = 10'd381;
assign feature_index_4[804] = 10'd247;
assign feature_index_4[805] = 10'd515;
assign feature_index_4[806] = 10'd0;
assign feature_index_4[807] = 10'd655;
assign feature_index_4[808] = 10'd156;
assign feature_index_4[809] = 10'd485;
assign feature_index_4[810] = 10'd401;
assign feature_index_4[811] = 10'd0;
assign feature_index_4[812] = 10'd0;
assign feature_index_4[813] = 10'd264;
assign feature_index_4[814] = 10'd265;
assign feature_index_4[815] = 10'd375;
assign feature_index_4[816] = 10'd515;
assign feature_index_4[817] = 10'd432;
assign feature_index_4[818] = 10'd430;
assign feature_index_4[819] = 10'd181;
assign feature_index_4[820] = 10'd628;
assign feature_index_4[821] = 10'd407;
assign feature_index_4[822] = 10'd377;
assign feature_index_4[823] = 10'd298;
assign feature_index_4[824] = 10'd239;
assign feature_index_4[825] = 10'd0;
assign feature_index_4[826] = 10'd205;
assign feature_index_4[827] = 10'd553;
assign feature_index_4[828] = 10'd382;
assign feature_index_4[829] = 10'd491;
assign feature_index_4[830] = 10'd426;
assign feature_index_4[831] = 10'd265;
assign feature_index_4[832] = 10'd332;
assign feature_index_4[833] = 10'd271;
assign feature_index_4[834] = 10'd570;
assign feature_index_4[835] = 10'd0;
assign feature_index_4[836] = 10'd149;
assign feature_index_4[837] = 10'd384;
assign feature_index_4[838] = 10'd295;
assign feature_index_4[839] = 10'd207;
assign feature_index_4[840] = 10'd0;
assign feature_index_4[841] = 10'd216;
assign feature_index_4[842] = 10'd0;
assign feature_index_4[843] = 10'd0;
assign feature_index_4[844] = 10'd600;
assign feature_index_4[845] = 10'd214;
assign feature_index_4[846] = 10'd0;
assign feature_index_4[847] = 10'd294;
assign feature_index_4[848] = 10'd347;
assign feature_index_4[849] = 10'd443;
assign feature_index_4[850] = 10'd649;
assign feature_index_4[851] = 10'd379;
assign feature_index_4[852] = 10'd543;
assign feature_index_4[853] = 10'd125;
assign feature_index_4[854] = 10'd380;
assign feature_index_4[855] = 10'd398;
assign feature_index_4[856] = 10'd99;
assign feature_index_4[857] = 10'd270;
assign feature_index_4[858] = 10'd468;
assign feature_index_4[859] = 10'd273;
assign feature_index_4[860] = 10'd680;
assign feature_index_4[861] = 10'd0;
assign feature_index_4[862] = 10'd288;
assign feature_index_4[863] = 10'd297;
assign feature_index_4[864] = 10'd0;
assign feature_index_4[865] = 10'd0;
assign feature_index_4[866] = 10'd0;
assign feature_index_4[867] = 10'd0;
assign feature_index_4[868] = 10'd0;
assign feature_index_4[869] = 10'd267;
assign feature_index_4[870] = 10'd0;
assign feature_index_4[871] = 10'd0;
assign feature_index_4[872] = 10'd0;
assign feature_index_4[873] = 10'd0;
assign feature_index_4[874] = 10'd0;
assign feature_index_4[875] = 10'd0;
assign feature_index_4[876] = 10'd0;
assign feature_index_4[877] = 10'd0;
assign feature_index_4[878] = 10'd0;
assign feature_index_4[879] = 10'd0;
assign feature_index_4[880] = 10'd0;
assign feature_index_4[881] = 10'd0;
assign feature_index_4[882] = 10'd0;
assign feature_index_4[883] = 10'd0;
assign feature_index_4[884] = 10'd0;
assign feature_index_4[885] = 10'd0;
assign feature_index_4[886] = 10'd0;
assign feature_index_4[887] = 10'd240;
assign feature_index_4[888] = 10'd0;
assign feature_index_4[889] = 10'd181;
assign feature_index_4[890] = 10'd0;
assign feature_index_4[891] = 10'd381;
assign feature_index_4[892] = 10'd410;
assign feature_index_4[893] = 10'd564;
assign feature_index_4[894] = 10'd276;
assign feature_index_4[895] = 10'd346;
assign feature_index_4[896] = 10'd482;
assign feature_index_4[897] = 10'd349;
assign feature_index_4[898] = 10'd160;
assign feature_index_4[899] = 10'd599;
assign feature_index_4[900] = 10'd71;
assign feature_index_4[901] = 10'd610;
assign feature_index_4[902] = 10'd260;
assign feature_index_4[903] = 10'd353;
assign feature_index_4[904] = 10'd487;
assign feature_index_4[905] = 10'd232;
assign feature_index_4[906] = 10'd624;
assign feature_index_4[907] = 10'd299;
assign feature_index_4[908] = 10'd632;
assign feature_index_4[909] = 10'd185;
assign feature_index_4[910] = 10'd130;
assign feature_index_4[911] = 10'd188;
assign feature_index_4[912] = 10'd0;
assign feature_index_4[913] = 10'd353;
assign feature_index_4[914] = 10'd320;
assign feature_index_4[915] = 10'd486;
assign feature_index_4[916] = 10'd264;
assign feature_index_4[917] = 10'd0;
assign feature_index_4[918] = 10'd348;
assign feature_index_4[919] = 10'd540;
assign feature_index_4[920] = 10'd0;
assign feature_index_4[921] = 10'd463;
assign feature_index_4[922] = 10'd459;
assign feature_index_4[923] = 10'd378;
assign feature_index_4[924] = 10'd602;
assign feature_index_4[925] = 10'd213;
assign feature_index_4[926] = 10'd400;
assign feature_index_4[927] = 10'd629;
assign feature_index_4[928] = 10'd300;
assign feature_index_4[929] = 10'd296;
assign feature_index_4[930] = 10'd181;
assign feature_index_4[931] = 10'd564;
assign feature_index_4[932] = 10'd93;
assign feature_index_4[933] = 10'd628;
assign feature_index_4[934] = 10'd626;
assign feature_index_4[935] = 10'd527;
assign feature_index_4[936] = 10'd433;
assign feature_index_4[937] = 10'd551;
assign feature_index_4[938] = 10'd0;
assign feature_index_4[939] = 10'd457;
assign feature_index_4[940] = 10'd267;
assign feature_index_4[941] = 10'd0;
assign feature_index_4[942] = 10'd495;
assign feature_index_4[943] = 10'd689;
assign feature_index_4[944] = 10'd215;
assign feature_index_4[945] = 10'd259;
assign feature_index_4[946] = 10'd405;
assign feature_index_4[947] = 10'd464;
assign feature_index_4[948] = 10'd0;
assign feature_index_4[949] = 10'd551;
assign feature_index_4[950] = 10'd192;
assign feature_index_4[951] = 10'd153;
assign feature_index_4[952] = 10'd0;
assign feature_index_4[953] = 10'd0;
assign feature_index_4[954] = 10'd211;
assign feature_index_4[955] = 10'd0;
assign feature_index_4[956] = 10'd0;
assign feature_index_4[957] = 10'd0;
assign feature_index_4[958] = 10'd233;
assign feature_index_4[959] = 10'd482;
assign feature_index_4[960] = 10'd98;
assign feature_index_4[961] = 10'd145;
assign feature_index_4[962] = 10'd626;
assign feature_index_4[963] = 10'd405;
assign feature_index_4[964] = 10'd463;
assign feature_index_4[965] = 10'd686;
assign feature_index_4[966] = 10'd0;
assign feature_index_4[967] = 10'd595;
assign feature_index_4[968] = 10'd410;
assign feature_index_4[969] = 10'd490;
assign feature_index_4[970] = 10'd434;
assign feature_index_4[971] = 10'd177;
assign feature_index_4[972] = 10'd636;
assign feature_index_4[973] = 10'd0;
assign feature_index_4[974] = 10'd0;
assign feature_index_4[975] = 10'd552;
assign feature_index_4[976] = 10'd515;
assign feature_index_4[977] = 10'd376;
assign feature_index_4[978] = 10'd368;
assign feature_index_4[979] = 10'd623;
assign feature_index_4[980] = 10'd436;
assign feature_index_4[981] = 10'd0;
assign feature_index_4[982] = 10'd240;
assign feature_index_4[983] = 10'd549;
assign feature_index_4[984] = 10'd510;
assign feature_index_4[985] = 10'd459;
assign feature_index_4[986] = 10'd512;
assign feature_index_4[987] = 10'd0;
assign feature_index_4[988] = 10'd0;
assign feature_index_4[989] = 10'd452;
assign feature_index_4[990] = 10'd536;
assign feature_index_4[991] = 10'd153;
assign feature_index_4[992] = 10'd457;
assign feature_index_4[993] = 10'd0;
assign feature_index_4[994] = 10'd683;
assign feature_index_4[995] = 10'd345;
assign feature_index_4[996] = 10'd0;
assign feature_index_4[997] = 10'd385;
assign feature_index_4[998] = 10'd0;
assign feature_index_4[999] = 10'd0;
assign feature_index_4[1000] = 10'd637;
assign feature_index_4[1001] = 10'd594;
assign feature_index_4[1002] = 10'd0;
assign feature_index_4[1003] = 10'd358;
assign feature_index_4[1004] = 10'd523;
assign feature_index_4[1005] = 10'd568;
assign feature_index_4[1006] = 10'd358;
assign feature_index_4[1007] = 10'd651;
assign feature_index_4[1008] = 10'd498;
assign feature_index_4[1009] = 10'd424;
assign feature_index_4[1010] = 10'd299;
assign feature_index_4[1011] = 10'd318;
assign feature_index_4[1012] = 10'd433;
assign feature_index_4[1013] = 10'd593;
assign feature_index_4[1014] = 10'd302;
assign feature_index_4[1015] = 10'd578;
assign feature_index_4[1016] = 10'd185;
assign feature_index_4[1017] = 10'd633;
assign feature_index_4[1018] = 10'd574;
assign feature_index_4[1019] = 10'd405;
assign feature_index_4[1020] = 10'd299;
assign feature_index_4[1021] = 10'd289;
assign feature_index_4[1022] = 10'd0;
assign feature_index_5[0] = 10'd378;
assign feature_index_5[1] = 10'd435;
assign feature_index_5[2] = 10'd410;
assign feature_index_5[3] = 10'd568;
assign feature_index_5[4] = 10'd268;
assign feature_index_5[5] = 10'd517;
assign feature_index_5[6] = 10'd487;
assign feature_index_5[7] = 10'd459;
assign feature_index_5[8] = 10'd516;
assign feature_index_5[9] = 10'd100;
assign feature_index_5[10] = 10'd431;
assign feature_index_5[11] = 10'd542;
assign feature_index_5[12] = 10'd318;
assign feature_index_5[13] = 10'd153;
assign feature_index_5[14] = 10'd654;
assign feature_index_5[15] = 10'd465;
assign feature_index_5[16] = 10'd653;
assign feature_index_5[17] = 10'd483;
assign feature_index_5[18] = 10'd414;
assign feature_index_5[19] = 10'd69;
assign feature_index_5[20] = 10'd298;
assign feature_index_5[21] = 10'd579;
assign feature_index_5[22] = 10'd569;
assign feature_index_5[23] = 10'd318;
assign feature_index_5[24] = 10'd290;
assign feature_index_5[25] = 10'd579;
assign feature_index_5[26] = 10'd441;
assign feature_index_5[27] = 10'd567;
assign feature_index_5[28] = 10'd295;
assign feature_index_5[29] = 10'd299;
assign feature_index_5[30] = 10'd456;
assign feature_index_5[31] = 10'd600;
assign feature_index_5[32] = 10'd483;
assign feature_index_5[33] = 10'd410;
assign feature_index_5[34] = 10'd384;
assign feature_index_5[35] = 10'd485;
assign feature_index_5[36] = 10'd301;
assign feature_index_5[37] = 10'd374;
assign feature_index_5[38] = 10'd125;
assign feature_index_5[39] = 10'd375;
assign feature_index_5[40] = 10'd564;
assign feature_index_5[41] = 10'd215;
assign feature_index_5[42] = 10'd374;
assign feature_index_5[43] = 10'd485;
assign feature_index_5[44] = 10'd691;
assign feature_index_5[45] = 10'd623;
assign feature_index_5[46] = 10'd271;
assign feature_index_5[47] = 10'd466;
assign feature_index_5[48] = 10'd157;
assign feature_index_5[49] = 10'd655;
assign feature_index_5[50] = 10'd470;
assign feature_index_5[51] = 10'd234;
assign feature_index_5[52] = 10'd385;
assign feature_index_5[53] = 10'd632;
assign feature_index_5[54] = 10'd327;
assign feature_index_5[55] = 10'd238;
assign feature_index_5[56] = 10'd592;
assign feature_index_5[57] = 10'd273;
assign feature_index_5[58] = 10'd322;
assign feature_index_5[59] = 10'd658;
assign feature_index_5[60] = 10'd598;
assign feature_index_5[61] = 10'd317;
assign feature_index_5[62] = 10'd349;
assign feature_index_5[63] = 10'd183;
assign feature_index_5[64] = 10'd324;
assign feature_index_5[65] = 10'd351;
assign feature_index_5[66] = 10'd302;
assign feature_index_5[67] = 10'd100;
assign feature_index_5[68] = 10'd543;
assign feature_index_5[69] = 10'd437;
assign feature_index_5[70] = 10'd376;
assign feature_index_5[71] = 10'd482;
assign feature_index_5[72] = 10'd352;
assign feature_index_5[73] = 10'd433;
assign feature_index_5[74] = 10'd459;
assign feature_index_5[75] = 10'd324;
assign feature_index_5[76] = 10'd440;
assign feature_index_5[77] = 10'd370;
assign feature_index_5[78] = 10'd269;
assign feature_index_5[79] = 10'd541;
assign feature_index_5[80] = 10'd299;
assign feature_index_5[81] = 10'd270;
assign feature_index_5[82] = 10'd0;
assign feature_index_5[83] = 10'd273;
assign feature_index_5[84] = 10'd291;
assign feature_index_5[85] = 10'd243;
assign feature_index_5[86] = 10'd595;
assign feature_index_5[87] = 10'd154;
assign feature_index_5[88] = 10'd540;
assign feature_index_5[89] = 10'd370;
assign feature_index_5[90] = 10'd343;
assign feature_index_5[91] = 10'd237;
assign feature_index_5[92] = 10'd516;
assign feature_index_5[93] = 10'd180;
assign feature_index_5[94] = 10'd294;
assign feature_index_5[95] = 10'd683;
assign feature_index_5[96] = 10'd219;
assign feature_index_5[97] = 10'd381;
assign feature_index_5[98] = 10'd484;
assign feature_index_5[99] = 10'd574;
assign feature_index_5[100] = 10'd292;
assign feature_index_5[101] = 10'd299;
assign feature_index_5[102] = 10'd567;
assign feature_index_5[103] = 10'd299;
assign feature_index_5[104] = 10'd526;
assign feature_index_5[105] = 10'd487;
assign feature_index_5[106] = 10'd245;
assign feature_index_5[107] = 10'd487;
assign feature_index_5[108] = 10'd544;
assign feature_index_5[109] = 10'd436;
assign feature_index_5[110] = 10'd216;
assign feature_index_5[111] = 10'd210;
assign feature_index_5[112] = 10'd497;
assign feature_index_5[113] = 10'd99;
assign feature_index_5[114] = 10'd163;
assign feature_index_5[115] = 10'd160;
assign feature_index_5[116] = 10'd428;
assign feature_index_5[117] = 10'd96;
assign feature_index_5[118] = 10'd151;
assign feature_index_5[119] = 10'd601;
assign feature_index_5[120] = 10'd153;
assign feature_index_5[121] = 10'd209;
assign feature_index_5[122] = 10'd596;
assign feature_index_5[123] = 10'd177;
assign feature_index_5[124] = 10'd156;
assign feature_index_5[125] = 10'd125;
assign feature_index_5[126] = 10'd379;
assign feature_index_5[127] = 10'd467;
assign feature_index_5[128] = 10'd538;
assign feature_index_5[129] = 10'd461;
assign feature_index_5[130] = 10'd453;
assign feature_index_5[131] = 10'd514;
assign feature_index_5[132] = 10'd316;
assign feature_index_5[133] = 10'd519;
assign feature_index_5[134] = 10'd510;
assign feature_index_5[135] = 10'd356;
assign feature_index_5[136] = 10'd563;
assign feature_index_5[137] = 10'd346;
assign feature_index_5[138] = 10'd656;
assign feature_index_5[139] = 10'd470;
assign feature_index_5[140] = 10'd188;
assign feature_index_5[141] = 10'd681;
assign feature_index_5[142] = 10'd515;
assign feature_index_5[143] = 10'd400;
assign feature_index_5[144] = 10'd403;
assign feature_index_5[145] = 10'd457;
assign feature_index_5[146] = 10'd291;
assign feature_index_5[147] = 10'd208;
assign feature_index_5[148] = 10'd298;
assign feature_index_5[149] = 10'd692;
assign feature_index_5[150] = 10'd347;
assign feature_index_5[151] = 10'd316;
assign feature_index_5[152] = 10'd174;
assign feature_index_5[153] = 10'd551;
assign feature_index_5[154] = 10'd186;
assign feature_index_5[155] = 10'd347;
assign feature_index_5[156] = 10'd229;
assign feature_index_5[157] = 10'd461;
assign feature_index_5[158] = 10'd461;
assign feature_index_5[159] = 10'd209;
assign feature_index_5[160] = 10'd398;
assign feature_index_5[161] = 10'd157;
assign feature_index_5[162] = 10'd597;
assign feature_index_5[163] = 10'd210;
assign feature_index_5[164] = 10'd494;
assign feature_index_5[165] = 10'd0;
assign feature_index_5[166] = 10'd0;
assign feature_index_5[167] = 10'd550;
assign feature_index_5[168] = 10'd318;
assign feature_index_5[169] = 10'd344;
assign feature_index_5[170] = 10'd162;
assign feature_index_5[171] = 10'd344;
assign feature_index_5[172] = 10'd0;
assign feature_index_5[173] = 10'd404;
assign feature_index_5[174] = 10'd292;
assign feature_index_5[175] = 10'd566;
assign feature_index_5[176] = 10'd321;
assign feature_index_5[177] = 10'd157;
assign feature_index_5[178] = 10'd428;
assign feature_index_5[179] = 10'd373;
assign feature_index_5[180] = 10'd210;
assign feature_index_5[181] = 10'd460;
assign feature_index_5[182] = 10'd183;
assign feature_index_5[183] = 10'd683;
assign feature_index_5[184] = 10'd376;
assign feature_index_5[185] = 10'd554;
assign feature_index_5[186] = 10'd488;
assign feature_index_5[187] = 10'd125;
assign feature_index_5[188] = 10'd632;
assign feature_index_5[189] = 10'd659;
assign feature_index_5[190] = 10'd383;
assign feature_index_5[191] = 10'd215;
assign feature_index_5[192] = 10'd513;
assign feature_index_5[193] = 10'd288;
assign feature_index_5[194] = 10'd430;
assign feature_index_5[195] = 10'd351;
assign feature_index_5[196] = 10'd520;
assign feature_index_5[197] = 10'd325;
assign feature_index_5[198] = 10'd497;
assign feature_index_5[199] = 10'd466;
assign feature_index_5[200] = 10'd180;
assign feature_index_5[201] = 10'd178;
assign feature_index_5[202] = 10'd373;
assign feature_index_5[203] = 10'd466;
assign feature_index_5[204] = 10'd380;
assign feature_index_5[205] = 10'd243;
assign feature_index_5[206] = 10'd239;
assign feature_index_5[207] = 10'd510;
assign feature_index_5[208] = 10'd297;
assign feature_index_5[209] = 10'd321;
assign feature_index_5[210] = 10'd359;
assign feature_index_5[211] = 10'd149;
assign feature_index_5[212] = 10'd689;
assign feature_index_5[213] = 10'd327;
assign feature_index_5[214] = 10'd184;
assign feature_index_5[215] = 10'd598;
assign feature_index_5[216] = 10'd185;
assign feature_index_5[217] = 10'd299;
assign feature_index_5[218] = 10'd581;
assign feature_index_5[219] = 10'd596;
assign feature_index_5[220] = 10'd458;
assign feature_index_5[221] = 10'd523;
assign feature_index_5[222] = 10'd359;
assign feature_index_5[223] = 10'd408;
assign feature_index_5[224] = 10'd321;
assign feature_index_5[225] = 10'd404;
assign feature_index_5[226] = 10'd228;
assign feature_index_5[227] = 10'd175;
assign feature_index_5[228] = 10'd426;
assign feature_index_5[229] = 10'd299;
assign feature_index_5[230] = 10'd462;
assign feature_index_5[231] = 10'd262;
assign feature_index_5[232] = 10'd651;
assign feature_index_5[233] = 10'd368;
assign feature_index_5[234] = 10'd631;
assign feature_index_5[235] = 10'd628;
assign feature_index_5[236] = 10'd0;
assign feature_index_5[237] = 10'd268;
assign feature_index_5[238] = 10'd191;
assign feature_index_5[239] = 10'd571;
assign feature_index_5[240] = 10'd575;
assign feature_index_5[241] = 10'd236;
assign feature_index_5[242] = 10'd489;
assign feature_index_5[243] = 10'd508;
assign feature_index_5[244] = 10'd188;
assign feature_index_5[245] = 10'd548;
assign feature_index_5[246] = 10'd291;
assign feature_index_5[247] = 10'd466;
assign feature_index_5[248] = 10'd610;
assign feature_index_5[249] = 10'd540;
assign feature_index_5[250] = 10'd272;
assign feature_index_5[251] = 10'd577;
assign feature_index_5[252] = 10'd437;
assign feature_index_5[253] = 10'd204;
assign feature_index_5[254] = 10'd274;
assign feature_index_5[255] = 10'd442;
assign feature_index_5[256] = 10'd655;
assign feature_index_5[257] = 10'd271;
assign feature_index_5[258] = 10'd244;
assign feature_index_5[259] = 10'd174;
assign feature_index_5[260] = 10'd495;
assign feature_index_5[261] = 10'd662;
assign feature_index_5[262] = 10'd269;
assign feature_index_5[263] = 10'd176;
assign feature_index_5[264] = 10'd517;
assign feature_index_5[265] = 10'd182;
assign feature_index_5[266] = 10'd154;
assign feature_index_5[267] = 10'd689;
assign feature_index_5[268] = 10'd210;
assign feature_index_5[269] = 10'd544;
assign feature_index_5[270] = 10'd185;
assign feature_index_5[271] = 10'd544;
assign feature_index_5[272] = 10'd324;
assign feature_index_5[273] = 10'd493;
assign feature_index_5[274] = 10'd0;
assign feature_index_5[275] = 10'd234;
assign feature_index_5[276] = 10'd711;
assign feature_index_5[277] = 10'd344;
assign feature_index_5[278] = 10'd347;
assign feature_index_5[279] = 10'd263;
assign feature_index_5[280] = 10'd295;
assign feature_index_5[281] = 10'd0;
assign feature_index_5[282] = 10'd658;
assign feature_index_5[283] = 10'd569;
assign feature_index_5[284] = 10'd548;
assign feature_index_5[285] = 10'd578;
assign feature_index_5[286] = 10'd377;
assign feature_index_5[287] = 10'd123;
assign feature_index_5[288] = 10'd535;
assign feature_index_5[289] = 10'd453;
assign feature_index_5[290] = 10'd207;
assign feature_index_5[291] = 10'd323;
assign feature_index_5[292] = 10'd429;
assign feature_index_5[293] = 10'd637;
assign feature_index_5[294] = 10'd401;
assign feature_index_5[295] = 10'd460;
assign feature_index_5[296] = 10'd351;
assign feature_index_5[297] = 10'd553;
assign feature_index_5[298] = 10'd351;
assign feature_index_5[299] = 10'd67;
assign feature_index_5[300] = 10'd655;
assign feature_index_5[301] = 10'd268;
assign feature_index_5[302] = 10'd489;
assign feature_index_5[303] = 10'd712;
assign feature_index_5[304] = 10'd426;
assign feature_index_5[305] = 10'd158;
assign feature_index_5[306] = 10'd0;
assign feature_index_5[307] = 10'd131;
assign feature_index_5[308] = 10'd124;
assign feature_index_5[309] = 10'd571;
assign feature_index_5[310] = 10'd552;
assign feature_index_5[311] = 10'd179;
assign feature_index_5[312] = 10'd399;
assign feature_index_5[313] = 10'd398;
assign feature_index_5[314] = 10'd604;
assign feature_index_5[315] = 10'd630;
assign feature_index_5[316] = 10'd467;
assign feature_index_5[317] = 10'd621;
assign feature_index_5[318] = 10'd0;
assign feature_index_5[319] = 10'd155;
assign feature_index_5[320] = 10'd598;
assign feature_index_5[321] = 10'd371;
assign feature_index_5[322] = 10'd182;
assign feature_index_5[323] = 10'd184;
assign feature_index_5[324] = 10'd541;
assign feature_index_5[325] = 10'd241;
assign feature_index_5[326] = 10'd455;
assign feature_index_5[327] = 10'd262;
assign feature_index_5[328] = 10'd294;
assign feature_index_5[329] = 10'd0;
assign feature_index_5[330] = 10'd0;
assign feature_index_5[331] = 10'd0;
assign feature_index_5[332] = 10'd0;
assign feature_index_5[333] = 10'd0;
assign feature_index_5[334] = 10'd0;
assign feature_index_5[335] = 10'd101;
assign feature_index_5[336] = 10'd623;
assign feature_index_5[337] = 10'd443;
assign feature_index_5[338] = 10'd0;
assign feature_index_5[339] = 10'd0;
assign feature_index_5[340] = 10'd567;
assign feature_index_5[341] = 10'd610;
assign feature_index_5[342] = 10'd342;
assign feature_index_5[343] = 10'd0;
assign feature_index_5[344] = 10'd0;
assign feature_index_5[345] = 10'd0;
assign feature_index_5[346] = 10'd0;
assign feature_index_5[347] = 10'd548;
assign feature_index_5[348] = 10'd412;
assign feature_index_5[349] = 10'd0;
assign feature_index_5[350] = 10'd349;
assign feature_index_5[351] = 10'd432;
assign feature_index_5[352] = 10'd455;
assign feature_index_5[353] = 10'd130;
assign feature_index_5[354] = 10'd482;
assign feature_index_5[355] = 10'd296;
assign feature_index_5[356] = 10'd324;
assign feature_index_5[357] = 10'd404;
assign feature_index_5[358] = 10'd131;
assign feature_index_5[359] = 10'd744;
assign feature_index_5[360] = 10'd574;
assign feature_index_5[361] = 10'd353;
assign feature_index_5[362] = 10'd572;
assign feature_index_5[363] = 10'd572;
assign feature_index_5[364] = 10'd156;
assign feature_index_5[365] = 10'd689;
assign feature_index_5[366] = 10'd412;
assign feature_index_5[367] = 10'd214;
assign feature_index_5[368] = 10'd545;
assign feature_index_5[369] = 10'd345;
assign feature_index_5[370] = 10'd379;
assign feature_index_5[371] = 10'd122;
assign feature_index_5[372] = 10'd631;
assign feature_index_5[373] = 10'd155;
assign feature_index_5[374] = 10'd539;
assign feature_index_5[375] = 10'd320;
assign feature_index_5[376] = 10'd354;
assign feature_index_5[377] = 10'd333;
assign feature_index_5[378] = 10'd216;
assign feature_index_5[379] = 10'd710;
assign feature_index_5[380] = 10'd657;
assign feature_index_5[381] = 10'd516;
assign feature_index_5[382] = 10'd460;
assign feature_index_5[383] = 10'd465;
assign feature_index_5[384] = 10'd151;
assign feature_index_5[385] = 10'd315;
assign feature_index_5[386] = 10'd353;
assign feature_index_5[387] = 10'd658;
assign feature_index_5[388] = 10'd152;
assign feature_index_5[389] = 10'd351;
assign feature_index_5[390] = 10'd650;
assign feature_index_5[391] = 10'd243;
assign feature_index_5[392] = 10'd217;
assign feature_index_5[393] = 10'd148;
assign feature_index_5[394] = 10'd623;
assign feature_index_5[395] = 10'd262;
assign feature_index_5[396] = 10'd269;
assign feature_index_5[397] = 10'd266;
assign feature_index_5[398] = 10'd654;
assign feature_index_5[399] = 10'd155;
assign feature_index_5[400] = 10'd600;
assign feature_index_5[401] = 10'd98;
assign feature_index_5[402] = 10'd292;
assign feature_index_5[403] = 10'd657;
assign feature_index_5[404] = 10'd493;
assign feature_index_5[405] = 10'd461;
assign feature_index_5[406] = 10'd634;
assign feature_index_5[407] = 10'd384;
assign feature_index_5[408] = 10'd515;
assign feature_index_5[409] = 10'd294;
assign feature_index_5[410] = 10'd438;
assign feature_index_5[411] = 10'd352;
assign feature_index_5[412] = 10'd358;
assign feature_index_5[413] = 10'd460;
assign feature_index_5[414] = 10'd303;
assign feature_index_5[415] = 10'd402;
assign feature_index_5[416] = 10'd178;
assign feature_index_5[417] = 10'd514;
assign feature_index_5[418] = 10'd275;
assign feature_index_5[419] = 10'd405;
assign feature_index_5[420] = 10'd655;
assign feature_index_5[421] = 10'd630;
assign feature_index_5[422] = 10'd0;
assign feature_index_5[423] = 10'd400;
assign feature_index_5[424] = 10'd472;
assign feature_index_5[425] = 10'd570;
assign feature_index_5[426] = 10'd572;
assign feature_index_5[427] = 10'd97;
assign feature_index_5[428] = 10'd691;
assign feature_index_5[429] = 10'd0;
assign feature_index_5[430] = 10'd286;
assign feature_index_5[431] = 10'd211;
assign feature_index_5[432] = 10'd353;
assign feature_index_5[433] = 10'd384;
assign feature_index_5[434] = 10'd272;
assign feature_index_5[435] = 10'd682;
assign feature_index_5[436] = 10'd326;
assign feature_index_5[437] = 10'd511;
assign feature_index_5[438] = 10'd465;
assign feature_index_5[439] = 10'd579;
assign feature_index_5[440] = 10'd386;
assign feature_index_5[441] = 10'd286;
assign feature_index_5[442] = 10'd102;
assign feature_index_5[443] = 10'd356;
assign feature_index_5[444] = 10'd571;
assign feature_index_5[445] = 10'd496;
assign feature_index_5[446] = 10'd570;
assign feature_index_5[447] = 10'd399;
assign feature_index_5[448] = 10'd283;
assign feature_index_5[449] = 10'd353;
assign feature_index_5[450] = 10'd490;
assign feature_index_5[451] = 10'd267;
assign feature_index_5[452] = 10'd159;
assign feature_index_5[453] = 10'd101;
assign feature_index_5[454] = 10'd427;
assign feature_index_5[455] = 10'd300;
assign feature_index_5[456] = 10'd441;
assign feature_index_5[457] = 10'd508;
assign feature_index_5[458] = 10'd0;
assign feature_index_5[459] = 10'd359;
assign feature_index_5[460] = 10'd208;
assign feature_index_5[461] = 10'd653;
assign feature_index_5[462] = 10'd459;
assign feature_index_5[463] = 10'd484;
assign feature_index_5[464] = 10'd356;
assign feature_index_5[465] = 10'd631;
assign feature_index_5[466] = 10'd161;
assign feature_index_5[467] = 10'd288;
assign feature_index_5[468] = 10'd0;
assign feature_index_5[469] = 10'd318;
assign feature_index_5[470] = 10'd467;
assign feature_index_5[471] = 10'd484;
assign feature_index_5[472] = 10'd123;
assign feature_index_5[473] = 10'd0;
assign feature_index_5[474] = 10'd0;
assign feature_index_5[475] = 10'd299;
assign feature_index_5[476] = 10'd135;
assign feature_index_5[477] = 10'd556;
assign feature_index_5[478] = 10'd296;
assign feature_index_5[479] = 10'd441;
assign feature_index_5[480] = 10'd538;
assign feature_index_5[481] = 10'd126;
assign feature_index_5[482] = 10'd203;
assign feature_index_5[483] = 10'd293;
assign feature_index_5[484] = 10'd404;
assign feature_index_5[485] = 10'd202;
assign feature_index_5[486] = 10'd635;
assign feature_index_5[487] = 10'd239;
assign feature_index_5[488] = 10'd386;
assign feature_index_5[489] = 10'd179;
assign feature_index_5[490] = 10'd630;
assign feature_index_5[491] = 10'd93;
assign feature_index_5[492] = 10'd688;
assign feature_index_5[493] = 10'd349;
assign feature_index_5[494] = 10'd347;
assign feature_index_5[495] = 10'd237;
assign feature_index_5[496] = 10'd542;
assign feature_index_5[497] = 10'd290;
assign feature_index_5[498] = 10'd567;
assign feature_index_5[499] = 10'd541;
assign feature_index_5[500] = 10'd256;
assign feature_index_5[501] = 10'd408;
assign feature_index_5[502] = 10'd425;
assign feature_index_5[503] = 10'd511;
assign feature_index_5[504] = 10'd191;
assign feature_index_5[505] = 10'd0;
assign feature_index_5[506] = 10'd341;
assign feature_index_5[507] = 10'd494;
assign feature_index_5[508] = 10'd442;
assign feature_index_5[509] = 10'd548;
assign feature_index_5[510] = 10'd512;
assign feature_index_5[511] = 10'd387;
assign feature_index_5[512] = 10'd341;
assign feature_index_5[513] = 10'd179;
assign feature_index_5[514] = 10'd351;
assign feature_index_5[515] = 10'd188;
assign feature_index_5[516] = 10'd542;
assign feature_index_5[517] = 10'd354;
assign feature_index_5[518] = 10'd321;
assign feature_index_5[519] = 10'd212;
assign feature_index_5[520] = 10'd571;
assign feature_index_5[521] = 10'd0;
assign feature_index_5[522] = 10'd0;
assign feature_index_5[523] = 10'd402;
assign feature_index_5[524] = 10'd512;
assign feature_index_5[525] = 10'd179;
assign feature_index_5[526] = 10'd0;
assign feature_index_5[527] = 10'd432;
assign feature_index_5[528] = 10'd150;
assign feature_index_5[529] = 10'd414;
assign feature_index_5[530] = 10'd567;
assign feature_index_5[531] = 10'd155;
assign feature_index_5[532] = 10'd402;
assign feature_index_5[533] = 10'd179;
assign feature_index_5[534] = 10'd152;
assign feature_index_5[535] = 10'd412;
assign feature_index_5[536] = 10'd601;
assign feature_index_5[537] = 10'd160;
assign feature_index_5[538] = 10'd654;
assign feature_index_5[539] = 10'd400;
assign feature_index_5[540] = 10'd124;
assign feature_index_5[541] = 10'd191;
assign feature_index_5[542] = 10'd652;
assign feature_index_5[543] = 10'd246;
assign feature_index_5[544] = 10'd128;
assign feature_index_5[545] = 10'd571;
assign feature_index_5[546] = 10'd457;
assign feature_index_5[547] = 10'd399;
assign feature_index_5[548] = 10'd0;
assign feature_index_5[549] = 10'd0;
assign feature_index_5[550] = 10'd0;
assign feature_index_5[551] = 10'd152;
assign feature_index_5[552] = 10'd601;
assign feature_index_5[553] = 10'd494;
assign feature_index_5[554] = 10'd409;
assign feature_index_5[555] = 10'd575;
assign feature_index_5[556] = 10'd574;
assign feature_index_5[557] = 10'd187;
assign feature_index_5[558] = 10'd230;
assign feature_index_5[559] = 10'd541;
assign feature_index_5[560] = 10'd0;
assign feature_index_5[561] = 10'd0;
assign feature_index_5[562] = 10'd0;
assign feature_index_5[563] = 10'd0;
assign feature_index_5[564] = 10'd0;
assign feature_index_5[565] = 10'd0;
assign feature_index_5[566] = 10'd0;
assign feature_index_5[567] = 10'd0;
assign feature_index_5[568] = 10'd0;
assign feature_index_5[569] = 10'd0;
assign feature_index_5[570] = 10'd484;
assign feature_index_5[571] = 10'd0;
assign feature_index_5[572] = 10'd0;
assign feature_index_5[573] = 10'd0;
assign feature_index_5[574] = 10'd0;
assign feature_index_5[575] = 10'd319;
assign feature_index_5[576] = 10'd289;
assign feature_index_5[577] = 10'd480;
assign feature_index_5[578] = 10'd265;
assign feature_index_5[579] = 10'd210;
assign feature_index_5[580] = 10'd370;
assign feature_index_5[581] = 10'd0;
assign feature_index_5[582] = 10'd0;
assign feature_index_5[583] = 10'd294;
assign feature_index_5[584] = 10'd0;
assign feature_index_5[585] = 10'd0;
assign feature_index_5[586] = 10'd272;
assign feature_index_5[587] = 10'd125;
assign feature_index_5[588] = 10'd0;
assign feature_index_5[589] = 10'd266;
assign feature_index_5[590] = 10'd269;
assign feature_index_5[591] = 10'd241;
assign feature_index_5[592] = 10'd188;
assign feature_index_5[593] = 10'd71;
assign feature_index_5[594] = 10'd686;
assign feature_index_5[595] = 10'd428;
assign feature_index_5[596] = 10'd0;
assign feature_index_5[597] = 10'd521;
assign feature_index_5[598] = 10'd130;
assign feature_index_5[599] = 10'd96;
assign feature_index_5[600] = 10'd0;
assign feature_index_5[601] = 10'd244;
assign feature_index_5[602] = 10'd0;
assign feature_index_5[603] = 10'd566;
assign feature_index_5[604] = 10'd491;
assign feature_index_5[605] = 10'd600;
assign feature_index_5[606] = 10'd387;
assign feature_index_5[607] = 10'd520;
assign feature_index_5[608] = 10'd0;
assign feature_index_5[609] = 10'd600;
assign feature_index_5[610] = 10'd441;
assign feature_index_5[611] = 10'd152;
assign feature_index_5[612] = 10'd73;
assign feature_index_5[613] = 10'd0;
assign feature_index_5[614] = 10'd0;
assign feature_index_5[615] = 10'd402;
assign feature_index_5[616] = 10'd576;
assign feature_index_5[617] = 10'd555;
assign feature_index_5[618] = 10'd547;
assign feature_index_5[619] = 10'd0;
assign feature_index_5[620] = 10'd498;
assign feature_index_5[621] = 10'd265;
assign feature_index_5[622] = 10'd206;
assign feature_index_5[623] = 10'd331;
assign feature_index_5[624] = 10'd192;
assign feature_index_5[625] = 10'd606;
assign feature_index_5[626] = 10'd488;
assign feature_index_5[627] = 10'd0;
assign feature_index_5[628] = 10'd303;
assign feature_index_5[629] = 10'd0;
assign feature_index_5[630] = 10'd0;
assign feature_index_5[631] = 10'd565;
assign feature_index_5[632] = 10'd624;
assign feature_index_5[633] = 10'd0;
assign feature_index_5[634] = 10'd0;
assign feature_index_5[635] = 10'd0;
assign feature_index_5[636] = 10'd319;
assign feature_index_5[637] = 10'd0;
assign feature_index_5[638] = 10'd0;
assign feature_index_5[639] = 10'd517;
assign feature_index_5[640] = 10'd345;
assign feature_index_5[641] = 10'd210;
assign feature_index_5[642] = 10'd372;
assign feature_index_5[643] = 10'd186;
assign feature_index_5[644] = 10'd443;
assign feature_index_5[645] = 10'd570;
assign feature_index_5[646] = 10'd572;
assign feature_index_5[647] = 10'd123;
assign feature_index_5[648] = 10'd325;
assign feature_index_5[649] = 10'd657;
assign feature_index_5[650] = 10'd301;
assign feature_index_5[651] = 10'd595;
assign feature_index_5[652] = 10'd469;
assign feature_index_5[653] = 10'd399;
assign feature_index_5[654] = 10'd581;
assign feature_index_5[655] = 10'd303;
assign feature_index_5[656] = 10'd0;
assign feature_index_5[657] = 10'd0;
assign feature_index_5[658] = 10'd460;
assign feature_index_5[659] = 10'd0;
assign feature_index_5[660] = 10'd0;
assign feature_index_5[661] = 10'd0;
assign feature_index_5[662] = 10'd0;
assign feature_index_5[663] = 10'd0;
assign feature_index_5[664] = 10'd0;
assign feature_index_5[665] = 10'd0;
assign feature_index_5[666] = 10'd0;
assign feature_index_5[667] = 10'd0;
assign feature_index_5[668] = 10'd0;
assign feature_index_5[669] = 10'd0;
assign feature_index_5[670] = 10'd0;
assign feature_index_5[671] = 10'd185;
assign feature_index_5[672] = 10'd184;
assign feature_index_5[673] = 10'd204;
assign feature_index_5[674] = 10'd346;
assign feature_index_5[675] = 10'd0;
assign feature_index_5[676] = 10'd0;
assign feature_index_5[677] = 10'd0;
assign feature_index_5[678] = 10'd0;
assign feature_index_5[679] = 10'd0;
assign feature_index_5[680] = 10'd0;
assign feature_index_5[681] = 10'd0;
assign feature_index_5[682] = 10'd0;
assign feature_index_5[683] = 10'd0;
assign feature_index_5[684] = 10'd0;
assign feature_index_5[685] = 10'd0;
assign feature_index_5[686] = 10'd0;
assign feature_index_5[687] = 10'd0;
assign feature_index_5[688] = 10'd0;
assign feature_index_5[689] = 10'd0;
assign feature_index_5[690] = 10'd0;
assign feature_index_5[691] = 10'd0;
assign feature_index_5[692] = 10'd0;
assign feature_index_5[693] = 10'd0;
assign feature_index_5[694] = 10'd0;
assign feature_index_5[695] = 10'd436;
assign feature_index_5[696] = 10'd0;
assign feature_index_5[697] = 10'd0;
assign feature_index_5[698] = 10'd0;
assign feature_index_5[699] = 10'd0;
assign feature_index_5[700] = 10'd0;
assign feature_index_5[701] = 10'd0;
assign feature_index_5[702] = 10'd467;
assign feature_index_5[703] = 10'd486;
assign feature_index_5[704] = 10'd410;
assign feature_index_5[705] = 10'd155;
assign feature_index_5[706] = 10'd273;
assign feature_index_5[707] = 10'd244;
assign feature_index_5[708] = 10'd541;
assign feature_index_5[709] = 10'd661;
assign feature_index_5[710] = 10'd650;
assign feature_index_5[711] = 10'd458;
assign feature_index_5[712] = 10'd372;
assign feature_index_5[713] = 10'd492;
assign feature_index_5[714] = 10'd327;
assign feature_index_5[715] = 10'd680;
assign feature_index_5[716] = 10'd484;
assign feature_index_5[717] = 10'd399;
assign feature_index_5[718] = 10'd218;
assign feature_index_5[719] = 10'd685;
assign feature_index_5[720] = 10'd0;
assign feature_index_5[721] = 10'd237;
assign feature_index_5[722] = 10'd401;
assign feature_index_5[723] = 10'd0;
assign feature_index_5[724] = 10'd328;
assign feature_index_5[725] = 10'd463;
assign feature_index_5[726] = 10'd541;
assign feature_index_5[727] = 10'd485;
assign feature_index_5[728] = 10'd666;
assign feature_index_5[729] = 10'd205;
assign feature_index_5[730] = 10'd345;
assign feature_index_5[731] = 10'd237;
assign feature_index_5[732] = 10'd271;
assign feature_index_5[733] = 10'd0;
assign feature_index_5[734] = 10'd523;
assign feature_index_5[735] = 10'd628;
assign feature_index_5[736] = 10'd294;
assign feature_index_5[737] = 10'd244;
assign feature_index_5[738] = 10'd601;
assign feature_index_5[739] = 10'd545;
assign feature_index_5[740] = 10'd324;
assign feature_index_5[741] = 10'd350;
assign feature_index_5[742] = 10'd288;
assign feature_index_5[743] = 10'd453;
assign feature_index_5[744] = 10'd293;
assign feature_index_5[745] = 10'd0;
assign feature_index_5[746] = 10'd372;
assign feature_index_5[747] = 10'd0;
assign feature_index_5[748] = 10'd0;
assign feature_index_5[749] = 10'd127;
assign feature_index_5[750] = 10'd579;
assign feature_index_5[751] = 10'd628;
assign feature_index_5[752] = 10'd485;
assign feature_index_5[753] = 10'd349;
assign feature_index_5[754] = 10'd0;
assign feature_index_5[755] = 10'd192;
assign feature_index_5[756] = 10'd0;
assign feature_index_5[757] = 10'd289;
assign feature_index_5[758] = 10'd178;
assign feature_index_5[759] = 10'd490;
assign feature_index_5[760] = 10'd0;
assign feature_index_5[761] = 10'd443;
assign feature_index_5[762] = 10'd684;
assign feature_index_5[763] = 10'd388;
assign feature_index_5[764] = 10'd380;
assign feature_index_5[765] = 10'd653;
assign feature_index_5[766] = 10'd402;
assign feature_index_5[767] = 10'd269;
assign feature_index_5[768] = 10'd627;
assign feature_index_5[769] = 10'd483;
assign feature_index_5[770] = 10'd464;
assign feature_index_5[771] = 10'd351;
assign feature_index_5[772] = 10'd369;
assign feature_index_5[773] = 10'd270;
assign feature_index_5[774] = 10'd496;
assign feature_index_5[775] = 10'd484;
assign feature_index_5[776] = 10'd178;
assign feature_index_5[777] = 10'd371;
assign feature_index_5[778] = 10'd346;
assign feature_index_5[779] = 10'd0;
assign feature_index_5[780] = 10'd265;
assign feature_index_5[781] = 10'd511;
assign feature_index_5[782] = 10'd463;
assign feature_index_5[783] = 10'd322;
assign feature_index_5[784] = 10'd493;
assign feature_index_5[785] = 10'd519;
assign feature_index_5[786] = 10'd414;
assign feature_index_5[787] = 10'd463;
assign feature_index_5[788] = 10'd594;
assign feature_index_5[789] = 10'd265;
assign feature_index_5[790] = 10'd513;
assign feature_index_5[791] = 10'd218;
assign feature_index_5[792] = 10'd425;
assign feature_index_5[793] = 10'd411;
assign feature_index_5[794] = 10'd152;
assign feature_index_5[795] = 10'd354;
assign feature_index_5[796] = 10'd353;
assign feature_index_5[797] = 10'd239;
assign feature_index_5[798] = 10'd382;
assign feature_index_5[799] = 10'd509;
assign feature_index_5[800] = 10'd576;
assign feature_index_5[801] = 10'd343;
assign feature_index_5[802] = 10'd610;
assign feature_index_5[803] = 10'd245;
assign feature_index_5[804] = 10'd437;
assign feature_index_5[805] = 10'd319;
assign feature_index_5[806] = 10'd457;
assign feature_index_5[807] = 10'd623;
assign feature_index_5[808] = 10'd515;
assign feature_index_5[809] = 10'd440;
assign feature_index_5[810] = 10'd608;
assign feature_index_5[811] = 10'd347;
assign feature_index_5[812] = 10'd432;
assign feature_index_5[813] = 10'd243;
assign feature_index_5[814] = 10'd357;
assign feature_index_5[815] = 10'd324;
assign feature_index_5[816] = 10'd656;
assign feature_index_5[817] = 10'd576;
assign feature_index_5[818] = 10'd269;
assign feature_index_5[819] = 10'd657;
assign feature_index_5[820] = 10'd383;
assign feature_index_5[821] = 10'd584;
assign feature_index_5[822] = 10'd564;
assign feature_index_5[823] = 10'd549;
assign feature_index_5[824] = 10'd582;
assign feature_index_5[825] = 10'd467;
assign feature_index_5[826] = 10'd609;
assign feature_index_5[827] = 10'd415;
assign feature_index_5[828] = 10'd555;
assign feature_index_5[829] = 10'd663;
assign feature_index_5[830] = 10'd0;
assign feature_index_5[831] = 10'd178;
assign feature_index_5[832] = 10'd550;
assign feature_index_5[833] = 10'd527;
assign feature_index_5[834] = 10'd0;
assign feature_index_5[835] = 10'd464;
assign feature_index_5[836] = 10'd536;
assign feature_index_5[837] = 10'd237;
assign feature_index_5[838] = 10'd651;
assign feature_index_5[839] = 10'd124;
assign feature_index_5[840] = 10'd576;
assign feature_index_5[841] = 10'd348;
assign feature_index_5[842] = 10'd680;
assign feature_index_5[843] = 10'd609;
assign feature_index_5[844] = 10'd540;
assign feature_index_5[845] = 10'd0;
assign feature_index_5[846] = 10'd0;
assign feature_index_5[847] = 10'd269;
assign feature_index_5[848] = 10'd484;
assign feature_index_5[849] = 10'd685;
assign feature_index_5[850] = 10'd331;
assign feature_index_5[851] = 10'd602;
assign feature_index_5[852] = 10'd387;
assign feature_index_5[853] = 10'd460;
assign feature_index_5[854] = 10'd316;
assign feature_index_5[855] = 10'd272;
assign feature_index_5[856] = 10'd0;
assign feature_index_5[857] = 10'd206;
assign feature_index_5[858] = 10'd0;
assign feature_index_5[859] = 10'd0;
assign feature_index_5[860] = 10'd0;
assign feature_index_5[861] = 10'd0;
assign feature_index_5[862] = 10'd0;
assign feature_index_5[863] = 10'd515;
assign feature_index_5[864] = 10'd634;
assign feature_index_5[865] = 10'd597;
assign feature_index_5[866] = 10'd569;
assign feature_index_5[867] = 10'd301;
assign feature_index_5[868] = 10'd271;
assign feature_index_5[869] = 10'd485;
assign feature_index_5[870] = 10'd629;
assign feature_index_5[871] = 10'd269;
assign feature_index_5[872] = 10'd513;
assign feature_index_5[873] = 10'd248;
assign feature_index_5[874] = 10'd398;
assign feature_index_5[875] = 10'd684;
assign feature_index_5[876] = 10'd600;
assign feature_index_5[877] = 10'd380;
assign feature_index_5[878] = 10'd317;
assign feature_index_5[879] = 10'd523;
assign feature_index_5[880] = 10'd0;
assign feature_index_5[881] = 10'd0;
assign feature_index_5[882] = 10'd105;
assign feature_index_5[883] = 10'd465;
assign feature_index_5[884] = 10'd546;
assign feature_index_5[885] = 10'd148;
assign feature_index_5[886] = 10'd540;
assign feature_index_5[887] = 10'd295;
assign feature_index_5[888] = 10'd406;
assign feature_index_5[889] = 10'd427;
assign feature_index_5[890] = 10'd311;
assign feature_index_5[891] = 10'd0;
assign feature_index_5[892] = 10'd182;
assign feature_index_5[893] = 10'd519;
assign feature_index_5[894] = 10'd0;
assign feature_index_5[895] = 10'd432;
assign feature_index_5[896] = 10'd338;
assign feature_index_5[897] = 10'd541;
assign feature_index_5[898] = 10'd405;
assign feature_index_5[899] = 10'd270;
assign feature_index_5[900] = 10'd184;
assign feature_index_5[901] = 10'd596;
assign feature_index_5[902] = 10'd266;
assign feature_index_5[903] = 10'd494;
assign feature_index_5[904] = 10'd233;
assign feature_index_5[905] = 10'd415;
assign feature_index_5[906] = 10'd245;
assign feature_index_5[907] = 10'd296;
assign feature_index_5[908] = 10'd0;
assign feature_index_5[909] = 10'd187;
assign feature_index_5[910] = 10'd260;
assign feature_index_5[911] = 10'd432;
assign feature_index_5[912] = 10'd346;
assign feature_index_5[913] = 10'd220;
assign feature_index_5[914] = 10'd206;
assign feature_index_5[915] = 10'd429;
assign feature_index_5[916] = 10'd0;
assign feature_index_5[917] = 10'd0;
assign feature_index_5[918] = 10'd0;
assign feature_index_5[919] = 10'd597;
assign feature_index_5[920] = 10'd0;
assign feature_index_5[921] = 10'd409;
assign feature_index_5[922] = 10'd582;
assign feature_index_5[923] = 10'd0;
assign feature_index_5[924] = 10'd432;
assign feature_index_5[925] = 10'd0;
assign feature_index_5[926] = 10'd0;
assign feature_index_5[927] = 10'd351;
assign feature_index_5[928] = 10'd291;
assign feature_index_5[929] = 10'd300;
assign feature_index_5[930] = 10'd514;
assign feature_index_5[931] = 10'd463;
assign feature_index_5[932] = 10'd658;
assign feature_index_5[933] = 10'd270;
assign feature_index_5[934] = 10'd348;
assign feature_index_5[935] = 10'd325;
assign feature_index_5[936] = 10'd469;
assign feature_index_5[937] = 10'd0;
assign feature_index_5[938] = 10'd0;
assign feature_index_5[939] = 10'd464;
assign feature_index_5[940] = 10'd568;
assign feature_index_5[941] = 10'd626;
assign feature_index_5[942] = 10'd541;
assign feature_index_5[943] = 10'd317;
assign feature_index_5[944] = 10'd349;
assign feature_index_5[945] = 10'd245;
assign feature_index_5[946] = 10'd599;
assign feature_index_5[947] = 10'd0;
assign feature_index_5[948] = 10'd0;
assign feature_index_5[949] = 10'd0;
assign feature_index_5[950] = 10'd0;
assign feature_index_5[951] = 10'd271;
assign feature_index_5[952] = 10'd350;
assign feature_index_5[953] = 10'd516;
assign feature_index_5[954] = 10'd0;
assign feature_index_5[955] = 10'd237;
assign feature_index_5[956] = 10'd203;
assign feature_index_5[957] = 10'd0;
assign feature_index_5[958] = 10'd267;
assign feature_index_5[959] = 10'd207;
assign feature_index_5[960] = 10'd324;
assign feature_index_5[961] = 10'd351;
assign feature_index_5[962] = 10'd153;
assign feature_index_5[963] = 10'd298;
assign feature_index_5[964] = 10'd343;
assign feature_index_5[965] = 10'd216;
assign feature_index_5[966] = 10'd268;
assign feature_index_5[967] = 10'd493;
assign feature_index_5[968] = 10'd270;
assign feature_index_5[969] = 10'd401;
assign feature_index_5[970] = 10'd598;
assign feature_index_5[971] = 10'd542;
assign feature_index_5[972] = 10'd371;
assign feature_index_5[973] = 10'd374;
assign feature_index_5[974] = 10'd145;
assign feature_index_5[975] = 10'd555;
assign feature_index_5[976] = 10'd711;
assign feature_index_5[977] = 10'd0;
assign feature_index_5[978] = 10'd571;
assign feature_index_5[979] = 10'd469;
assign feature_index_5[980] = 10'd261;
assign feature_index_5[981] = 10'd659;
assign feature_index_5[982] = 10'd628;
assign feature_index_5[983] = 10'd497;
assign feature_index_5[984] = 10'd0;
assign feature_index_5[985] = 10'd656;
assign feature_index_5[986] = 10'd522;
assign feature_index_5[987] = 10'd574;
assign feature_index_5[988] = 10'd526;
assign feature_index_5[989] = 10'd679;
assign feature_index_5[990] = 10'd442;
assign feature_index_5[991] = 10'd324;
assign feature_index_5[992] = 10'd486;
assign feature_index_5[993] = 10'd320;
assign feature_index_5[994] = 10'd292;
assign feature_index_5[995] = 10'd657;
assign feature_index_5[996] = 10'd401;
assign feature_index_5[997] = 10'd575;
assign feature_index_5[998] = 10'd429;
assign feature_index_5[999] = 10'd660;
assign feature_index_5[1000] = 10'd686;
assign feature_index_5[1001] = 10'd649;
assign feature_index_5[1002] = 10'd148;
assign feature_index_5[1003] = 10'd205;
assign feature_index_5[1004] = 10'd515;
assign feature_index_5[1005] = 10'd347;
assign feature_index_5[1006] = 10'd0;
assign feature_index_5[1007] = 10'd542;
assign feature_index_5[1008] = 10'd630;
assign feature_index_5[1009] = 10'd373;
assign feature_index_5[1010] = 10'd329;
assign feature_index_5[1011] = 10'd0;
assign feature_index_5[1012] = 10'd0;
assign feature_index_5[1013] = 10'd0;
assign feature_index_5[1014] = 10'd584;
assign feature_index_5[1015] = 10'd606;
assign feature_index_5[1016] = 10'd0;
assign feature_index_5[1017] = 10'd0;
assign feature_index_5[1018] = 10'd0;
assign feature_index_5[1019] = 10'd183;
assign feature_index_5[1020] = 10'd573;
assign feature_index_5[1021] = 10'd156;
assign feature_index_5[1022] = 10'd452;
assign feature_index_6[0] = 10'd539;
assign feature_index_6[1] = 10'd261;
assign feature_index_6[2] = 10'd317;
assign feature_index_6[3] = 10'd347;
assign feature_index_6[4] = 10'd459;
assign feature_index_6[5] = 10'd153;
assign feature_index_6[6] = 10'd405;
assign feature_index_6[7] = 10'd437;
assign feature_index_6[8] = 10'd711;
assign feature_index_6[9] = 10'd402;
assign feature_index_6[10] = 10'd240;
assign feature_index_6[11] = 10'd320;
assign feature_index_6[12] = 10'd629;
assign feature_index_6[13] = 10'd628;
assign feature_index_6[14] = 10'd513;
assign feature_index_6[15] = 10'd577;
assign feature_index_6[16] = 10'd179;
assign feature_index_6[17] = 10'd178;
assign feature_index_6[18] = 10'd213;
assign feature_index_6[19] = 10'd153;
assign feature_index_6[20] = 10'd239;
assign feature_index_6[21] = 10'd96;
assign feature_index_6[22] = 10'd400;
assign feature_index_6[23] = 10'd491;
assign feature_index_6[24] = 10'd654;
assign feature_index_6[25] = 10'd314;
assign feature_index_6[26] = 10'd459;
assign feature_index_6[27] = 10'd269;
assign feature_index_6[28] = 10'd456;
assign feature_index_6[29] = 10'd329;
assign feature_index_6[30] = 10'd299;
assign feature_index_6[31] = 10'd235;
assign feature_index_6[32] = 10'd488;
assign feature_index_6[33] = 10'd264;
assign feature_index_6[34] = 10'd153;
assign feature_index_6[35] = 10'd551;
assign feature_index_6[36] = 10'd625;
assign feature_index_6[37] = 10'd737;
assign feature_index_6[38] = 10'd408;
assign feature_index_6[39] = 10'd156;
assign feature_index_6[40] = 10'd352;
assign feature_index_6[41] = 10'd552;
assign feature_index_6[42] = 10'd633;
assign feature_index_6[43] = 10'd350;
assign feature_index_6[44] = 10'd215;
assign feature_index_6[45] = 10'd345;
assign feature_index_6[46] = 10'd569;
assign feature_index_6[47] = 10'd650;
assign feature_index_6[48] = 10'd237;
assign feature_index_6[49] = 10'd522;
assign feature_index_6[50] = 10'd373;
assign feature_index_6[51] = 10'd375;
assign feature_index_6[52] = 10'd577;
assign feature_index_6[53] = 10'd323;
assign feature_index_6[54] = 10'd265;
assign feature_index_6[55] = 10'd435;
assign feature_index_6[56] = 10'd441;
assign feature_index_6[57] = 10'd324;
assign feature_index_6[58] = 10'd432;
assign feature_index_6[59] = 10'd325;
assign feature_index_6[60] = 10'd398;
assign feature_index_6[61] = 10'd100;
assign feature_index_6[62] = 10'd187;
assign feature_index_6[63] = 10'd205;
assign feature_index_6[64] = 10'd214;
assign feature_index_6[65] = 10'd345;
assign feature_index_6[66] = 10'd294;
assign feature_index_6[67] = 10'd597;
assign feature_index_6[68] = 10'd206;
assign feature_index_6[69] = 10'd523;
assign feature_index_6[70] = 10'd541;
assign feature_index_6[71] = 10'd624;
assign feature_index_6[72] = 10'd595;
assign feature_index_6[73] = 10'd290;
assign feature_index_6[74] = 10'd236;
assign feature_index_6[75] = 10'd461;
assign feature_index_6[76] = 10'd459;
assign feature_index_6[77] = 10'd173;
assign feature_index_6[78] = 10'd574;
assign feature_index_6[79] = 10'd377;
assign feature_index_6[80] = 10'd347;
assign feature_index_6[81] = 10'd378;
assign feature_index_6[82] = 10'd489;
assign feature_index_6[83] = 10'd156;
assign feature_index_6[84] = 10'd376;
assign feature_index_6[85] = 10'd622;
assign feature_index_6[86] = 10'd188;
assign feature_index_6[87] = 10'd456;
assign feature_index_6[88] = 10'd429;
assign feature_index_6[89] = 10'd273;
assign feature_index_6[90] = 10'd185;
assign feature_index_6[91] = 10'd343;
assign feature_index_6[92] = 10'd182;
assign feature_index_6[93] = 10'd176;
assign feature_index_6[94] = 10'd542;
assign feature_index_6[95] = 10'd313;
assign feature_index_6[96] = 10'd269;
assign feature_index_6[97] = 10'd286;
assign feature_index_6[98] = 10'd602;
assign feature_index_6[99] = 10'd411;
assign feature_index_6[100] = 10'd462;
assign feature_index_6[101] = 10'd512;
assign feature_index_6[102] = 10'd184;
assign feature_index_6[103] = 10'd488;
assign feature_index_6[104] = 10'd679;
assign feature_index_6[105] = 10'd379;
assign feature_index_6[106] = 10'd453;
assign feature_index_6[107] = 10'd408;
assign feature_index_6[108] = 10'd291;
assign feature_index_6[109] = 10'd321;
assign feature_index_6[110] = 10'd435;
assign feature_index_6[111] = 10'd437;
assign feature_index_6[112] = 10'd215;
assign feature_index_6[113] = 10'd416;
assign feature_index_6[114] = 10'd354;
assign feature_index_6[115] = 10'd369;
assign feature_index_6[116] = 10'd330;
assign feature_index_6[117] = 10'd490;
assign feature_index_6[118] = 10'd212;
assign feature_index_6[119] = 10'd358;
assign feature_index_6[120] = 10'd457;
assign feature_index_6[121] = 10'd523;
assign feature_index_6[122] = 10'd295;
assign feature_index_6[123] = 10'd244;
assign feature_index_6[124] = 10'd209;
assign feature_index_6[125] = 10'd516;
assign feature_index_6[126] = 10'd400;
assign feature_index_6[127] = 10'd406;
assign feature_index_6[128] = 10'd455;
assign feature_index_6[129] = 10'd176;
assign feature_index_6[130] = 10'd292;
assign feature_index_6[131] = 10'd203;
assign feature_index_6[132] = 10'd523;
assign feature_index_6[133] = 10'd542;
assign feature_index_6[134] = 10'd610;
assign feature_index_6[135] = 10'd428;
assign feature_index_6[136] = 10'd294;
assign feature_index_6[137] = 10'd160;
assign feature_index_6[138] = 10'd550;
assign feature_index_6[139] = 10'd399;
assign feature_index_6[140] = 10'd635;
assign feature_index_6[141] = 10'd490;
assign feature_index_6[142] = 10'd348;
assign feature_index_6[143] = 10'd345;
assign feature_index_6[144] = 10'd569;
assign feature_index_6[145] = 10'd659;
assign feature_index_6[146] = 10'd426;
assign feature_index_6[147] = 10'd260;
assign feature_index_6[148] = 10'd69;
assign feature_index_6[149] = 10'd513;
assign feature_index_6[150] = 10'd269;
assign feature_index_6[151] = 10'd405;
assign feature_index_6[152] = 10'd188;
assign feature_index_6[153] = 10'd406;
assign feature_index_6[154] = 10'd240;
assign feature_index_6[155] = 10'd327;
assign feature_index_6[156] = 10'd0;
assign feature_index_6[157] = 10'd292;
assign feature_index_6[158] = 10'd432;
assign feature_index_6[159] = 10'd513;
assign feature_index_6[160] = 10'd317;
assign feature_index_6[161] = 10'd397;
assign feature_index_6[162] = 10'd460;
assign feature_index_6[163] = 10'd435;
assign feature_index_6[164] = 10'd322;
assign feature_index_6[165] = 10'd405;
assign feature_index_6[166] = 10'd349;
assign feature_index_6[167] = 10'd182;
assign feature_index_6[168] = 10'd461;
assign feature_index_6[169] = 10'd213;
assign feature_index_6[170] = 10'd454;
assign feature_index_6[171] = 10'd263;
assign feature_index_6[172] = 10'd298;
assign feature_index_6[173] = 10'd489;
assign feature_index_6[174] = 10'd300;
assign feature_index_6[175] = 10'd182;
assign feature_index_6[176] = 10'd182;
assign feature_index_6[177] = 10'd271;
assign feature_index_6[178] = 10'd572;
assign feature_index_6[179] = 10'd271;
assign feature_index_6[180] = 10'd573;
assign feature_index_6[181] = 10'd0;
assign feature_index_6[182] = 10'd0;
assign feature_index_6[183] = 10'd348;
assign feature_index_6[184] = 10'd456;
assign feature_index_6[185] = 10'd243;
assign feature_index_6[186] = 10'd214;
assign feature_index_6[187] = 10'd356;
assign feature_index_6[188] = 10'd684;
assign feature_index_6[189] = 10'd344;
assign feature_index_6[190] = 10'd524;
assign feature_index_6[191] = 10'd486;
assign feature_index_6[192] = 10'd353;
assign feature_index_6[193] = 10'd208;
assign feature_index_6[194] = 10'd488;
assign feature_index_6[195] = 10'd551;
assign feature_index_6[196] = 10'd387;
assign feature_index_6[197] = 10'd285;
assign feature_index_6[198] = 10'd655;
assign feature_index_6[199] = 10'd458;
assign feature_index_6[200] = 10'd462;
assign feature_index_6[201] = 10'd384;
assign feature_index_6[202] = 10'd299;
assign feature_index_6[203] = 10'd682;
assign feature_index_6[204] = 10'd353;
assign feature_index_6[205] = 10'd355;
assign feature_index_6[206] = 10'd220;
assign feature_index_6[207] = 10'd492;
assign feature_index_6[208] = 10'd517;
assign feature_index_6[209] = 10'd440;
assign feature_index_6[210] = 10'd0;
assign feature_index_6[211] = 10'd275;
assign feature_index_6[212] = 10'd607;
assign feature_index_6[213] = 10'd416;
assign feature_index_6[214] = 10'd354;
assign feature_index_6[215] = 10'd370;
assign feature_index_6[216] = 10'd150;
assign feature_index_6[217] = 10'd399;
assign feature_index_6[218] = 10'd296;
assign feature_index_6[219] = 10'd571;
assign feature_index_6[220] = 10'd580;
assign feature_index_6[221] = 10'd346;
assign feature_index_6[222] = 10'd513;
assign feature_index_6[223] = 10'd380;
assign feature_index_6[224] = 10'd415;
assign feature_index_6[225] = 10'd547;
assign feature_index_6[226] = 10'd239;
assign feature_index_6[227] = 10'd425;
assign feature_index_6[228] = 10'd381;
assign feature_index_6[229] = 10'd415;
assign feature_index_6[230] = 10'd360;
assign feature_index_6[231] = 10'd387;
assign feature_index_6[232] = 10'd510;
assign feature_index_6[233] = 10'd266;
assign feature_index_6[234] = 10'd242;
assign feature_index_6[235] = 10'd400;
assign feature_index_6[236] = 10'd434;
assign feature_index_6[237] = 10'd601;
assign feature_index_6[238] = 10'd414;
assign feature_index_6[239] = 10'd326;
assign feature_index_6[240] = 10'd303;
assign feature_index_6[241] = 10'd274;
assign feature_index_6[242] = 10'd571;
assign feature_index_6[243] = 10'd411;
assign feature_index_6[244] = 10'd484;
assign feature_index_6[245] = 10'd127;
assign feature_index_6[246] = 10'd177;
assign feature_index_6[247] = 10'd544;
assign feature_index_6[248] = 10'd407;
assign feature_index_6[249] = 10'd135;
assign feature_index_6[250] = 10'd573;
assign feature_index_6[251] = 10'd265;
assign feature_index_6[252] = 10'd427;
assign feature_index_6[253] = 10'd246;
assign feature_index_6[254] = 10'd408;
assign feature_index_6[255] = 10'd131;
assign feature_index_6[256] = 10'd291;
assign feature_index_6[257] = 10'd634;
assign feature_index_6[258] = 10'd246;
assign feature_index_6[259] = 10'd320;
assign feature_index_6[260] = 10'd288;
assign feature_index_6[261] = 10'd152;
assign feature_index_6[262] = 10'd406;
assign feature_index_6[263] = 10'd439;
assign feature_index_6[264] = 10'd483;
assign feature_index_6[265] = 10'd129;
assign feature_index_6[266] = 10'd603;
assign feature_index_6[267] = 10'd404;
assign feature_index_6[268] = 10'd385;
assign feature_index_6[269] = 10'd552;
assign feature_index_6[270] = 10'd0;
assign feature_index_6[271] = 10'd349;
assign feature_index_6[272] = 10'd570;
assign feature_index_6[273] = 10'd681;
assign feature_index_6[274] = 10'd487;
assign feature_index_6[275] = 10'd156;
assign feature_index_6[276] = 10'd508;
assign feature_index_6[277] = 10'd555;
assign feature_index_6[278] = 10'd631;
assign feature_index_6[279] = 10'd578;
assign feature_index_6[280] = 10'd204;
assign feature_index_6[281] = 10'd349;
assign feature_index_6[282] = 10'd657;
assign feature_index_6[283] = 10'd346;
assign feature_index_6[284] = 10'd377;
assign feature_index_6[285] = 10'd349;
assign feature_index_6[286] = 10'd176;
assign feature_index_6[287] = 10'd572;
assign feature_index_6[288] = 10'd399;
assign feature_index_6[289] = 10'd571;
assign feature_index_6[290] = 10'd516;
assign feature_index_6[291] = 10'd575;
assign feature_index_6[292] = 10'd434;
assign feature_index_6[293] = 10'd190;
assign feature_index_6[294] = 10'd408;
assign feature_index_6[295] = 10'd287;
assign feature_index_6[296] = 10'd461;
assign feature_index_6[297] = 10'd210;
assign feature_index_6[298] = 10'd0;
assign feature_index_6[299] = 10'd296;
assign feature_index_6[300] = 10'd463;
assign feature_index_6[301] = 10'd262;
assign feature_index_6[302] = 10'd262;
assign feature_index_6[303] = 10'd295;
assign feature_index_6[304] = 10'd204;
assign feature_index_6[305] = 10'd400;
assign feature_index_6[306] = 10'd0;
assign feature_index_6[307] = 10'd484;
assign feature_index_6[308] = 10'd654;
assign feature_index_6[309] = 10'd0;
assign feature_index_6[310] = 10'd0;
assign feature_index_6[311] = 10'd217;
assign feature_index_6[312] = 10'd183;
assign feature_index_6[313] = 10'd0;
assign feature_index_6[314] = 10'd0;
assign feature_index_6[315] = 10'd488;
assign feature_index_6[316] = 10'd521;
assign feature_index_6[317] = 10'd379;
assign feature_index_6[318] = 10'd628;
assign feature_index_6[319] = 10'd525;
assign feature_index_6[320] = 10'd182;
assign feature_index_6[321] = 10'd183;
assign feature_index_6[322] = 10'd325;
assign feature_index_6[323] = 10'd518;
assign feature_index_6[324] = 10'd463;
assign feature_index_6[325] = 10'd302;
assign feature_index_6[326] = 10'd0;
assign feature_index_6[327] = 10'd381;
assign feature_index_6[328] = 10'd300;
assign feature_index_6[329] = 10'd356;
assign feature_index_6[330] = 10'd516;
assign feature_index_6[331] = 10'd291;
assign feature_index_6[332] = 10'd323;
assign feature_index_6[333] = 10'd414;
assign feature_index_6[334] = 10'd320;
assign feature_index_6[335] = 10'd124;
assign feature_index_6[336] = 10'd488;
assign feature_index_6[337] = 10'd375;
assign feature_index_6[338] = 10'd600;
assign feature_index_6[339] = 10'd602;
assign feature_index_6[340] = 10'd342;
assign feature_index_6[341] = 10'd326;
assign feature_index_6[342] = 10'd429;
assign feature_index_6[343] = 10'd466;
assign feature_index_6[344] = 10'd431;
assign feature_index_6[345] = 10'd513;
assign feature_index_6[346] = 10'd455;
assign feature_index_6[347] = 10'd457;
assign feature_index_6[348] = 10'd522;
assign feature_index_6[349] = 10'd489;
assign feature_index_6[350] = 10'd432;
assign feature_index_6[351] = 10'd441;
assign feature_index_6[352] = 10'd486;
assign feature_index_6[353] = 10'd499;
assign feature_index_6[354] = 10'd98;
assign feature_index_6[355] = 10'd517;
assign feature_index_6[356] = 10'd717;
assign feature_index_6[357] = 10'd568;
assign feature_index_6[358] = 10'd655;
assign feature_index_6[359] = 10'd239;
assign feature_index_6[360] = 10'd156;
assign feature_index_6[361] = 10'd0;
assign feature_index_6[362] = 10'd0;
assign feature_index_6[363] = 10'd0;
assign feature_index_6[364] = 10'd0;
assign feature_index_6[365] = 10'd0;
assign feature_index_6[366] = 10'd0;
assign feature_index_6[367] = 10'd153;
assign feature_index_6[368] = 10'd550;
assign feature_index_6[369] = 10'd573;
assign feature_index_6[370] = 10'd469;
assign feature_index_6[371] = 10'd266;
assign feature_index_6[372] = 10'd381;
assign feature_index_6[373] = 10'd378;
assign feature_index_6[374] = 10'd571;
assign feature_index_6[375] = 10'd238;
assign feature_index_6[376] = 10'd438;
assign feature_index_6[377] = 10'd266;
assign feature_index_6[378] = 10'd518;
assign feature_index_6[379] = 10'd209;
assign feature_index_6[380] = 10'd576;
assign feature_index_6[381] = 10'd435;
assign feature_index_6[382] = 10'd434;
assign feature_index_6[383] = 10'd324;
assign feature_index_6[384] = 10'd371;
assign feature_index_6[385] = 10'd410;
assign feature_index_6[386] = 10'd181;
assign feature_index_6[387] = 10'd188;
assign feature_index_6[388] = 10'd592;
assign feature_index_6[389] = 10'd485;
assign feature_index_6[390] = 10'd211;
assign feature_index_6[391] = 10'd100;
assign feature_index_6[392] = 10'd466;
assign feature_index_6[393] = 10'd353;
assign feature_index_6[394] = 10'd201;
assign feature_index_6[395] = 10'd655;
assign feature_index_6[396] = 10'd267;
assign feature_index_6[397] = 10'd687;
assign feature_index_6[398] = 10'd405;
assign feature_index_6[399] = 10'd414;
assign feature_index_6[400] = 10'd157;
assign feature_index_6[401] = 10'd624;
assign feature_index_6[402] = 10'd302;
assign feature_index_6[403] = 10'd330;
assign feature_index_6[404] = 10'd216;
assign feature_index_6[405] = 10'd217;
assign feature_index_6[406] = 10'd183;
assign feature_index_6[407] = 10'd258;
assign feature_index_6[408] = 10'd219;
assign feature_index_6[409] = 10'd402;
assign feature_index_6[410] = 10'd494;
assign feature_index_6[411] = 10'd413;
assign feature_index_6[412] = 10'd400;
assign feature_index_6[413] = 10'd428;
assign feature_index_6[414] = 10'd300;
assign feature_index_6[415] = 10'd440;
assign feature_index_6[416] = 10'd460;
assign feature_index_6[417] = 10'd315;
assign feature_index_6[418] = 10'd163;
assign feature_index_6[419] = 10'd608;
assign feature_index_6[420] = 10'd491;
assign feature_index_6[421] = 10'd0;
assign feature_index_6[422] = 10'd0;
assign feature_index_6[423] = 10'd567;
assign feature_index_6[424] = 10'd0;
assign feature_index_6[425] = 10'd296;
assign feature_index_6[426] = 10'd285;
assign feature_index_6[427] = 10'd0;
assign feature_index_6[428] = 10'd0;
assign feature_index_6[429] = 10'd463;
assign feature_index_6[430] = 10'd357;
assign feature_index_6[431] = 10'd150;
assign feature_index_6[432] = 10'd434;
assign feature_index_6[433] = 10'd163;
assign feature_index_6[434] = 10'd94;
assign feature_index_6[435] = 10'd458;
assign feature_index_6[436] = 10'd443;
assign feature_index_6[437] = 10'd598;
assign feature_index_6[438] = 10'd124;
assign feature_index_6[439] = 10'd378;
assign feature_index_6[440] = 10'd457;
assign feature_index_6[441] = 10'd523;
assign feature_index_6[442] = 10'd410;
assign feature_index_6[443] = 10'd657;
assign feature_index_6[444] = 10'd215;
assign feature_index_6[445] = 10'd319;
assign feature_index_6[446] = 10'd608;
assign feature_index_6[447] = 10'd278;
assign feature_index_6[448] = 10'd294;
assign feature_index_6[449] = 10'd515;
assign feature_index_6[450] = 10'd217;
assign feature_index_6[451] = 10'd457;
assign feature_index_6[452] = 10'd592;
assign feature_index_6[453] = 10'd624;
assign feature_index_6[454] = 10'd654;
assign feature_index_6[455] = 10'd209;
assign feature_index_6[456] = 10'd213;
assign feature_index_6[457] = 10'd0;
assign feature_index_6[458] = 10'd0;
assign feature_index_6[459] = 10'd461;
assign feature_index_6[460] = 10'd163;
assign feature_index_6[461] = 10'd406;
assign feature_index_6[462] = 10'd319;
assign feature_index_6[463] = 10'd427;
assign feature_index_6[464] = 10'd409;
assign feature_index_6[465] = 10'd0;
assign feature_index_6[466] = 10'd584;
assign feature_index_6[467] = 10'd98;
assign feature_index_6[468] = 10'd218;
assign feature_index_6[469] = 10'd372;
assign feature_index_6[470] = 10'd207;
assign feature_index_6[471] = 10'd370;
assign feature_index_6[472] = 10'd473;
assign feature_index_6[473] = 10'd624;
assign feature_index_6[474] = 10'd712;
assign feature_index_6[475] = 10'd0;
assign feature_index_6[476] = 10'd127;
assign feature_index_6[477] = 10'd461;
assign feature_index_6[478] = 10'd524;
assign feature_index_6[479] = 10'd121;
assign feature_index_6[480] = 10'd379;
assign feature_index_6[481] = 10'd0;
assign feature_index_6[482] = 10'd0;
assign feature_index_6[483] = 10'd264;
assign feature_index_6[484] = 10'd157;
assign feature_index_6[485] = 10'd653;
assign feature_index_6[486] = 10'd517;
assign feature_index_6[487] = 10'd188;
assign feature_index_6[488] = 10'd493;
assign feature_index_6[489] = 10'd349;
assign feature_index_6[490] = 10'd374;
assign feature_index_6[491] = 10'd430;
assign feature_index_6[492] = 10'd489;
assign feature_index_6[493] = 10'd385;
assign feature_index_6[494] = 10'd0;
assign feature_index_6[495] = 10'd131;
assign feature_index_6[496] = 10'd583;
assign feature_index_6[497] = 10'd345;
assign feature_index_6[498] = 10'd191;
assign feature_index_6[499] = 10'd181;
assign feature_index_6[500] = 10'd0;
assign feature_index_6[501] = 10'd295;
assign feature_index_6[502] = 10'd243;
assign feature_index_6[503] = 10'd442;
assign feature_index_6[504] = 10'd570;
assign feature_index_6[505] = 10'd211;
assign feature_index_6[506] = 10'd369;
assign feature_index_6[507] = 10'd656;
assign feature_index_6[508] = 10'd582;
assign feature_index_6[509] = 10'd495;
assign feature_index_6[510] = 10'd659;
assign feature_index_6[511] = 10'd436;
assign feature_index_6[512] = 10'd524;
assign feature_index_6[513] = 10'd663;
assign feature_index_6[514] = 10'd469;
assign feature_index_6[515] = 10'd229;
assign feature_index_6[516] = 10'd685;
assign feature_index_6[517] = 10'd686;
assign feature_index_6[518] = 10'd0;
assign feature_index_6[519] = 10'd289;
assign feature_index_6[520] = 10'd157;
assign feature_index_6[521] = 10'd313;
assign feature_index_6[522] = 10'd0;
assign feature_index_6[523] = 10'd372;
assign feature_index_6[524] = 10'd543;
assign feature_index_6[525] = 10'd271;
assign feature_index_6[526] = 10'd604;
assign feature_index_6[527] = 10'd324;
assign feature_index_6[528] = 10'd187;
assign feature_index_6[529] = 10'd381;
assign feature_index_6[530] = 10'd627;
assign feature_index_6[531] = 10'd382;
assign feature_index_6[532] = 10'd325;
assign feature_index_6[533] = 10'd273;
assign feature_index_6[534] = 10'd407;
assign feature_index_6[535] = 10'd344;
assign feature_index_6[536] = 10'd346;
assign feature_index_6[537] = 10'd441;
assign feature_index_6[538] = 10'd244;
assign feature_index_6[539] = 10'd626;
assign feature_index_6[540] = 10'd456;
assign feature_index_6[541] = 10'd0;
assign feature_index_6[542] = 10'd0;
assign feature_index_6[543] = 10'd543;
assign feature_index_6[544] = 10'd655;
assign feature_index_6[545] = 10'd566;
assign feature_index_6[546] = 10'd372;
assign feature_index_6[547] = 10'd513;
assign feature_index_6[548] = 10'd268;
assign feature_index_6[549] = 10'd515;
assign feature_index_6[550] = 10'd324;
assign feature_index_6[551] = 10'd318;
assign feature_index_6[552] = 10'd657;
assign feature_index_6[553] = 10'd182;
assign feature_index_6[554] = 10'd544;
assign feature_index_6[555] = 10'd535;
assign feature_index_6[556] = 10'd0;
assign feature_index_6[557] = 10'd404;
assign feature_index_6[558] = 10'd0;
assign feature_index_6[559] = 10'd604;
assign feature_index_6[560] = 10'd546;
assign feature_index_6[561] = 10'd0;
assign feature_index_6[562] = 10'd233;
assign feature_index_6[563] = 10'd552;
assign feature_index_6[564] = 10'd712;
assign feature_index_6[565] = 10'd218;
assign feature_index_6[566] = 10'd314;
assign feature_index_6[567] = 10'd344;
assign feature_index_6[568] = 10'd542;
assign feature_index_6[569] = 10'd606;
assign feature_index_6[570] = 10'd629;
assign feature_index_6[571] = 10'd572;
assign feature_index_6[572] = 10'd245;
assign feature_index_6[573] = 10'd515;
assign feature_index_6[574] = 10'd626;
assign feature_index_6[575] = 10'd353;
assign feature_index_6[576] = 10'd522;
assign feature_index_6[577] = 10'd239;
assign feature_index_6[578] = 10'd267;
assign feature_index_6[579] = 10'd353;
assign feature_index_6[580] = 10'd351;
assign feature_index_6[581] = 10'd292;
assign feature_index_6[582] = 10'd657;
assign feature_index_6[583] = 10'd599;
assign feature_index_6[584] = 10'd213;
assign feature_index_6[585] = 10'd150;
assign feature_index_6[586] = 10'd208;
assign feature_index_6[587] = 10'd513;
assign feature_index_6[588] = 10'd555;
assign feature_index_6[589] = 10'd292;
assign feature_index_6[590] = 10'd564;
assign feature_index_6[591] = 10'd473;
assign feature_index_6[592] = 10'd400;
assign feature_index_6[593] = 10'd344;
assign feature_index_6[594] = 10'd631;
assign feature_index_6[595] = 10'd183;
assign feature_index_6[596] = 10'd327;
assign feature_index_6[597] = 10'd0;
assign feature_index_6[598] = 10'd0;
assign feature_index_6[599] = 10'd235;
assign feature_index_6[600] = 10'd349;
assign feature_index_6[601] = 10'd267;
assign feature_index_6[602] = 10'd286;
assign feature_index_6[603] = 10'd189;
assign feature_index_6[604] = 10'd328;
assign feature_index_6[605] = 10'd528;
assign feature_index_6[606] = 10'd466;
assign feature_index_6[607] = 10'd300;
assign feature_index_6[608] = 10'd204;
assign feature_index_6[609] = 10'd437;
assign feature_index_6[610] = 10'd0;
assign feature_index_6[611] = 10'd515;
assign feature_index_6[612] = 10'd240;
assign feature_index_6[613] = 10'd0;
assign feature_index_6[614] = 10'd0;
assign feature_index_6[615] = 10'd0;
assign feature_index_6[616] = 10'd0;
assign feature_index_6[617] = 10'd0;
assign feature_index_6[618] = 10'd0;
assign feature_index_6[619] = 10'd0;
assign feature_index_6[620] = 10'd0;
assign feature_index_6[621] = 10'd0;
assign feature_index_6[622] = 10'd0;
assign feature_index_6[623] = 10'd179;
assign feature_index_6[624] = 10'd355;
assign feature_index_6[625] = 10'd324;
assign feature_index_6[626] = 10'd217;
assign feature_index_6[627] = 10'd0;
assign feature_index_6[628] = 10'd0;
assign feature_index_6[629] = 10'd0;
assign feature_index_6[630] = 10'd0;
assign feature_index_6[631] = 10'd0;
assign feature_index_6[632] = 10'd301;
assign feature_index_6[633] = 10'd242;
assign feature_index_6[634] = 10'd301;
assign feature_index_6[635] = 10'd457;
assign feature_index_6[636] = 10'd378;
assign feature_index_6[637] = 10'd462;
assign feature_index_6[638] = 10'd248;
assign feature_index_6[639] = 10'd555;
assign feature_index_6[640] = 10'd510;
assign feature_index_6[641] = 10'd121;
assign feature_index_6[642] = 10'd554;
assign feature_index_6[643] = 10'd524;
assign feature_index_6[644] = 10'd232;
assign feature_index_6[645] = 10'd461;
assign feature_index_6[646] = 10'd329;
assign feature_index_6[647] = 10'd427;
assign feature_index_6[648] = 10'd513;
assign feature_index_6[649] = 10'd0;
assign feature_index_6[650] = 10'd682;
assign feature_index_6[651] = 10'd325;
assign feature_index_6[652] = 10'd0;
assign feature_index_6[653] = 10'd0;
assign feature_index_6[654] = 10'd0;
assign feature_index_6[655] = 10'd375;
assign feature_index_6[656] = 10'd482;
assign feature_index_6[657] = 10'd628;
assign feature_index_6[658] = 10'd376;
assign feature_index_6[659] = 10'd202;
assign feature_index_6[660] = 10'd248;
assign feature_index_6[661] = 10'd188;
assign feature_index_6[662] = 10'd426;
assign feature_index_6[663] = 10'd650;
assign feature_index_6[664] = 10'd202;
assign feature_index_6[665] = 10'd176;
assign feature_index_6[666] = 10'd485;
assign feature_index_6[667] = 10'd468;
assign feature_index_6[668] = 10'd185;
assign feature_index_6[669] = 10'd431;
assign feature_index_6[670] = 10'd469;
assign feature_index_6[671] = 10'd399;
assign feature_index_6[672] = 10'd624;
assign feature_index_6[673] = 10'd211;
assign feature_index_6[674] = 10'd403;
assign feature_index_6[675] = 10'd627;
assign feature_index_6[676] = 10'd318;
assign feature_index_6[677] = 10'd626;
assign feature_index_6[678] = 10'd400;
assign feature_index_6[679] = 10'd297;
assign feature_index_6[680] = 10'd484;
assign feature_index_6[681] = 10'd596;
assign feature_index_6[682] = 10'd0;
assign feature_index_6[683] = 10'd155;
assign feature_index_6[684] = 10'd272;
assign feature_index_6[685] = 10'd0;
assign feature_index_6[686] = 10'd596;
assign feature_index_6[687] = 10'd627;
assign feature_index_6[688] = 10'd243;
assign feature_index_6[689] = 10'd465;
assign feature_index_6[690] = 10'd409;
assign feature_index_6[691] = 10'd289;
assign feature_index_6[692] = 10'd0;
assign feature_index_6[693] = 10'd403;
assign feature_index_6[694] = 10'd601;
assign feature_index_6[695] = 10'd151;
assign feature_index_6[696] = 10'd377;
assign feature_index_6[697] = 10'd484;
assign feature_index_6[698] = 10'd554;
assign feature_index_6[699] = 10'd299;
assign feature_index_6[700] = 10'd191;
assign feature_index_6[701] = 10'd468;
assign feature_index_6[702] = 10'd597;
assign feature_index_6[703] = 10'd271;
assign feature_index_6[704] = 10'd465;
assign feature_index_6[705] = 10'd271;
assign feature_index_6[706] = 10'd566;
assign feature_index_6[707] = 10'd322;
assign feature_index_6[708] = 10'd299;
assign feature_index_6[709] = 10'd301;
assign feature_index_6[710] = 10'd516;
assign feature_index_6[711] = 10'd498;
assign feature_index_6[712] = 10'd184;
assign feature_index_6[713] = 10'd659;
assign feature_index_6[714] = 10'd0;
assign feature_index_6[715] = 10'd600;
assign feature_index_6[716] = 10'd580;
assign feature_index_6[717] = 10'd713;
assign feature_index_6[718] = 10'd546;
assign feature_index_6[719] = 10'd567;
assign feature_index_6[720] = 10'd376;
assign feature_index_6[721] = 10'd0;
assign feature_index_6[722] = 10'd0;
assign feature_index_6[723] = 10'd0;
assign feature_index_6[724] = 10'd0;
assign feature_index_6[725] = 10'd0;
assign feature_index_6[726] = 10'd0;
assign feature_index_6[727] = 10'd0;
assign feature_index_6[728] = 10'd0;
assign feature_index_6[729] = 10'd0;
assign feature_index_6[730] = 10'd0;
assign feature_index_6[731] = 10'd0;
assign feature_index_6[732] = 10'd0;
assign feature_index_6[733] = 10'd0;
assign feature_index_6[734] = 10'd0;
assign feature_index_6[735] = 10'd579;
assign feature_index_6[736] = 10'd581;
assign feature_index_6[737] = 10'd296;
assign feature_index_6[738] = 10'd515;
assign feature_index_6[739] = 10'd370;
assign feature_index_6[740] = 10'd570;
assign feature_index_6[741] = 10'd208;
assign feature_index_6[742] = 10'd580;
assign feature_index_6[743] = 10'd745;
assign feature_index_6[744] = 10'd654;
assign feature_index_6[745] = 10'd465;
assign feature_index_6[746] = 10'd266;
assign feature_index_6[747] = 10'd321;
assign feature_index_6[748] = 10'd627;
assign feature_index_6[749] = 10'd409;
assign feature_index_6[750] = 10'd379;
assign feature_index_6[751] = 10'd208;
assign feature_index_6[752] = 10'd409;
assign feature_index_6[753] = 10'd265;
assign feature_index_6[754] = 10'd178;
assign feature_index_6[755] = 10'd181;
assign feature_index_6[756] = 10'd369;
assign feature_index_6[757] = 10'd689;
assign feature_index_6[758] = 10'd442;
assign feature_index_6[759] = 10'd0;
assign feature_index_6[760] = 10'd0;
assign feature_index_6[761] = 10'd500;
assign feature_index_6[762] = 10'd369;
assign feature_index_6[763] = 10'd434;
assign feature_index_6[764] = 10'd287;
assign feature_index_6[765] = 10'd183;
assign feature_index_6[766] = 10'd689;
assign feature_index_6[767] = 10'd493;
assign feature_index_6[768] = 10'd359;
assign feature_index_6[769] = 10'd580;
assign feature_index_6[770] = 10'd324;
assign feature_index_6[771] = 10'd438;
assign feature_index_6[772] = 10'd433;
assign feature_index_6[773] = 10'd230;
assign feature_index_6[774] = 10'd412;
assign feature_index_6[775] = 10'd651;
assign feature_index_6[776] = 10'd0;
assign feature_index_6[777] = 10'd0;
assign feature_index_6[778] = 10'd0;
assign feature_index_6[779] = 10'd0;
assign feature_index_6[780] = 10'd631;
assign feature_index_6[781] = 10'd704;
assign feature_index_6[782] = 10'd356;
assign feature_index_6[783] = 10'd427;
assign feature_index_6[784] = 10'd182;
assign feature_index_6[785] = 10'd343;
assign feature_index_6[786] = 10'd0;
assign feature_index_6[787] = 10'd343;
assign feature_index_6[788] = 10'd636;
assign feature_index_6[789] = 10'd185;
assign feature_index_6[790] = 10'd376;
assign feature_index_6[791] = 10'd487;
assign feature_index_6[792] = 10'd297;
assign feature_index_6[793] = 10'd596;
assign feature_index_6[794] = 10'd547;
assign feature_index_6[795] = 10'd377;
assign feature_index_6[796] = 10'd383;
assign feature_index_6[797] = 10'd623;
assign feature_index_6[798] = 10'd321;
assign feature_index_6[799] = 10'd663;
assign feature_index_6[800] = 10'd0;
assign feature_index_6[801] = 10'd322;
assign feature_index_6[802] = 10'd347;
assign feature_index_6[803] = 10'd319;
assign feature_index_6[804] = 10'd497;
assign feature_index_6[805] = 10'd576;
assign feature_index_6[806] = 10'd572;
assign feature_index_6[807] = 10'd246;
assign feature_index_6[808] = 10'd358;
assign feature_index_6[809] = 10'd244;
assign feature_index_6[810] = 10'd375;
assign feature_index_6[811] = 10'd499;
assign feature_index_6[812] = 10'd104;
assign feature_index_6[813] = 10'd268;
assign feature_index_6[814] = 10'd101;
assign feature_index_6[815] = 10'd601;
assign feature_index_6[816] = 10'd229;
assign feature_index_6[817] = 10'd513;
assign feature_index_6[818] = 10'd356;
assign feature_index_6[819] = 10'd404;
assign feature_index_6[820] = 10'd246;
assign feature_index_6[821] = 10'd635;
assign feature_index_6[822] = 10'd405;
assign feature_index_6[823] = 10'd152;
assign feature_index_6[824] = 10'd0;
assign feature_index_6[825] = 10'd485;
assign feature_index_6[826] = 10'd380;
assign feature_index_6[827] = 10'd459;
assign feature_index_6[828] = 10'd266;
assign feature_index_6[829] = 10'd386;
assign feature_index_6[830] = 10'd351;
assign feature_index_6[831] = 10'd408;
assign feature_index_6[832] = 10'd454;
assign feature_index_6[833] = 10'd607;
assign feature_index_6[834] = 10'd0;
assign feature_index_6[835] = 10'd600;
assign feature_index_6[836] = 10'd0;
assign feature_index_6[837] = 10'd316;
assign feature_index_6[838] = 10'd351;
assign feature_index_6[839] = 10'd320;
assign feature_index_6[840] = 10'd0;
assign feature_index_6[841] = 10'd514;
assign feature_index_6[842] = 10'd101;
assign feature_index_6[843] = 10'd0;
assign feature_index_6[844] = 10'd0;
assign feature_index_6[845] = 10'd0;
assign feature_index_6[846] = 10'd0;
assign feature_index_6[847] = 10'd0;
assign feature_index_6[848] = 10'd432;
assign feature_index_6[849] = 10'd0;
assign feature_index_6[850] = 10'd0;
assign feature_index_6[851] = 10'd0;
assign feature_index_6[852] = 10'd0;
assign feature_index_6[853] = 10'd0;
assign feature_index_6[854] = 10'd0;
assign feature_index_6[855] = 10'd0;
assign feature_index_6[856] = 10'd0;
assign feature_index_6[857] = 10'd0;
assign feature_index_6[858] = 10'd0;
assign feature_index_6[859] = 10'd0;
assign feature_index_6[860] = 10'd0;
assign feature_index_6[861] = 10'd0;
assign feature_index_6[862] = 10'd547;
assign feature_index_6[863] = 10'd272;
assign feature_index_6[864] = 10'd350;
assign feature_index_6[865] = 10'd488;
assign feature_index_6[866] = 10'd0;
assign feature_index_6[867] = 10'd514;
assign feature_index_6[868] = 10'd654;
assign feature_index_6[869] = 10'd457;
assign feature_index_6[870] = 10'd0;
assign feature_index_6[871] = 10'd331;
assign feature_index_6[872] = 10'd668;
assign feature_index_6[873] = 10'd434;
assign feature_index_6[874] = 10'd382;
assign feature_index_6[875] = 10'd433;
assign feature_index_6[876] = 10'd591;
assign feature_index_6[877] = 10'd243;
assign feature_index_6[878] = 10'd463;
assign feature_index_6[879] = 10'd684;
assign feature_index_6[880] = 10'd437;
assign feature_index_6[881] = 10'd429;
assign feature_index_6[882] = 10'd341;
assign feature_index_6[883] = 10'd485;
assign feature_index_6[884] = 10'd548;
assign feature_index_6[885] = 10'd246;
assign feature_index_6[886] = 10'd241;
assign feature_index_6[887] = 10'd272;
assign feature_index_6[888] = 10'd324;
assign feature_index_6[889] = 10'd262;
assign feature_index_6[890] = 10'd540;
assign feature_index_6[891] = 10'd456;
assign feature_index_6[892] = 10'd385;
assign feature_index_6[893] = 10'd469;
assign feature_index_6[894] = 10'd212;
assign feature_index_6[895] = 10'd611;
assign feature_index_6[896] = 10'd0;
assign feature_index_6[897] = 10'd0;
assign feature_index_6[898] = 10'd0;
assign feature_index_6[899] = 10'd492;
assign feature_index_6[900] = 10'd442;
assign feature_index_6[901] = 10'd456;
assign feature_index_6[902] = 10'd179;
assign feature_index_6[903] = 10'd575;
assign feature_index_6[904] = 10'd519;
assign feature_index_6[905] = 10'd384;
assign feature_index_6[906] = 10'd211;
assign feature_index_6[907] = 10'd571;
assign feature_index_6[908] = 10'd412;
assign feature_index_6[909] = 10'd651;
assign feature_index_6[910] = 10'd623;
assign feature_index_6[911] = 10'd410;
assign feature_index_6[912] = 10'd525;
assign feature_index_6[913] = 10'd357;
assign feature_index_6[914] = 10'd440;
assign feature_index_6[915] = 10'd0;
assign feature_index_6[916] = 10'd0;
assign feature_index_6[917] = 10'd0;
assign feature_index_6[918] = 10'd0;
assign feature_index_6[919] = 10'd716;
assign feature_index_6[920] = 10'd570;
assign feature_index_6[921] = 10'd508;
assign feature_index_6[922] = 10'd0;
assign feature_index_6[923] = 10'd461;
assign feature_index_6[924] = 10'd385;
assign feature_index_6[925] = 10'd407;
assign feature_index_6[926] = 10'd0;
assign feature_index_6[927] = 10'd518;
assign feature_index_6[928] = 10'd408;
assign feature_index_6[929] = 10'd146;
assign feature_index_6[930] = 10'd412;
assign feature_index_6[931] = 10'd0;
assign feature_index_6[932] = 10'd0;
assign feature_index_6[933] = 10'd262;
assign feature_index_6[934] = 10'd662;
assign feature_index_6[935] = 10'd269;
assign feature_index_6[936] = 10'd520;
assign feature_index_6[937] = 10'd123;
assign feature_index_6[938] = 10'd347;
assign feature_index_6[939] = 10'd0;
assign feature_index_6[940] = 10'd374;
assign feature_index_6[941] = 10'd232;
assign feature_index_6[942] = 10'd497;
assign feature_index_6[943] = 10'd145;
assign feature_index_6[944] = 10'd638;
assign feature_index_6[945] = 10'd483;
assign feature_index_6[946] = 10'd315;
assign feature_index_6[947] = 10'd269;
assign feature_index_6[948] = 10'd583;
assign feature_index_6[949] = 10'd372;
assign feature_index_6[950] = 10'd0;
assign feature_index_6[951] = 10'd0;
assign feature_index_6[952] = 10'd0;
assign feature_index_6[953] = 10'd485;
assign feature_index_6[954] = 10'd242;
assign feature_index_6[955] = 10'd104;
assign feature_index_6[956] = 10'd152;
assign feature_index_6[957] = 10'd489;
assign feature_index_6[958] = 10'd371;
assign feature_index_6[959] = 10'd78;
assign feature_index_6[960] = 10'd494;
assign feature_index_6[961] = 10'd294;
assign feature_index_6[962] = 10'd465;
assign feature_index_6[963] = 10'd0;
assign feature_index_6[964] = 10'd0;
assign feature_index_6[965] = 10'd0;
assign feature_index_6[966] = 10'd0;
assign feature_index_6[967] = 10'd101;
assign feature_index_6[968] = 10'd358;
assign feature_index_6[969] = 10'd0;
assign feature_index_6[970] = 10'd299;
assign feature_index_6[971] = 10'd625;
assign feature_index_6[972] = 10'd621;
assign feature_index_6[973] = 10'd428;
assign feature_index_6[974] = 10'd463;
assign feature_index_6[975] = 10'd518;
assign feature_index_6[976] = 10'd717;
assign feature_index_6[977] = 10'd486;
assign feature_index_6[978] = 10'd428;
assign feature_index_6[979] = 10'd459;
assign feature_index_6[980] = 10'd0;
assign feature_index_6[981] = 10'd578;
assign feature_index_6[982] = 10'd187;
assign feature_index_6[983] = 10'd574;
assign feature_index_6[984] = 10'd380;
assign feature_index_6[985] = 10'd520;
assign feature_index_6[986] = 10'd316;
assign feature_index_6[987] = 10'd399;
assign feature_index_6[988] = 10'd106;
assign feature_index_6[989] = 10'd0;
assign feature_index_6[990] = 10'd0;
assign feature_index_6[991] = 10'd433;
assign feature_index_6[992] = 10'd661;
assign feature_index_6[993] = 10'd549;
assign feature_index_6[994] = 10'd268;
assign feature_index_6[995] = 10'd0;
assign feature_index_6[996] = 10'd433;
assign feature_index_6[997] = 10'd383;
assign feature_index_6[998] = 10'd384;
assign feature_index_6[999] = 10'd627;
assign feature_index_6[1000] = 10'd0;
assign feature_index_6[1001] = 10'd0;
assign feature_index_6[1002] = 10'd0;
assign feature_index_6[1003] = 10'd0;
assign feature_index_6[1004] = 10'd0;
assign feature_index_6[1005] = 10'd241;
assign feature_index_6[1006] = 10'd489;
assign feature_index_6[1007] = 10'd209;
assign feature_index_6[1008] = 10'd348;
assign feature_index_6[1009] = 10'd461;
assign feature_index_6[1010] = 10'd354;
assign feature_index_6[1011] = 10'd353;
assign feature_index_6[1012] = 10'd355;
assign feature_index_6[1013] = 10'd717;
assign feature_index_6[1014] = 10'd325;
assign feature_index_6[1015] = 10'd236;
assign feature_index_6[1016] = 10'd320;
assign feature_index_6[1017] = 10'd652;
assign feature_index_6[1018] = 10'd322;
assign feature_index_6[1019] = 10'd469;
assign feature_index_6[1020] = 10'd602;
assign feature_index_6[1021] = 10'd175;
assign feature_index_6[1022] = 10'd441;
assign feature_index_7[0] = 10'd461;
assign feature_index_7[1] = 10'd539;
assign feature_index_7[2] = 10'd347;
assign feature_index_7[3] = 10'd155;
assign feature_index_7[4] = 10'd442;
assign feature_index_7[5] = 10'd458;
assign feature_index_7[6] = 10'd103;
assign feature_index_7[7] = 10'd514;
assign feature_index_7[8] = 10'd428;
assign feature_index_7[9] = 10'd372;
assign feature_index_7[10] = 10'd343;
assign feature_index_7[11] = 10'd409;
assign feature_index_7[12] = 10'd540;
assign feature_index_7[13] = 10'd377;
assign feature_index_7[14] = 10'd211;
assign feature_index_7[15] = 10'd375;
assign feature_index_7[16] = 10'd96;
assign feature_index_7[17] = 10'd263;
assign feature_index_7[18] = 10'd406;
assign feature_index_7[19] = 10'd456;
assign feature_index_7[20] = 10'd350;
assign feature_index_7[21] = 10'd377;
assign feature_index_7[22] = 10'd352;
assign feature_index_7[23] = 10'd521;
assign feature_index_7[24] = 10'd710;
assign feature_index_7[25] = 10'd210;
assign feature_index_7[26] = 10'd656;
assign feature_index_7[27] = 10'd437;
assign feature_index_7[28] = 10'd100;
assign feature_index_7[29] = 10'd99;
assign feature_index_7[30] = 10'd378;
assign feature_index_7[31] = 10'd379;
assign feature_index_7[32] = 10'd622;
assign feature_index_7[33] = 10'd215;
assign feature_index_7[34] = 10'd158;
assign feature_index_7[35] = 10'd654;
assign feature_index_7[36] = 10'd268;
assign feature_index_7[37] = 10'd630;
assign feature_index_7[38] = 10'd288;
assign feature_index_7[39] = 10'd631;
assign feature_index_7[40] = 10'd346;
assign feature_index_7[41] = 10'd356;
assign feature_index_7[42] = 10'd456;
assign feature_index_7[43] = 10'd245;
assign feature_index_7[44] = 10'd274;
assign feature_index_7[45] = 10'd597;
assign feature_index_7[46] = 10'd296;
assign feature_index_7[47] = 10'd289;
assign feature_index_7[48] = 10'd373;
assign feature_index_7[49] = 10'd579;
assign feature_index_7[50] = 10'd430;
assign feature_index_7[51] = 10'd153;
assign feature_index_7[52] = 10'd262;
assign feature_index_7[53] = 10'd154;
assign feature_index_7[54] = 10'd153;
assign feature_index_7[55] = 10'd523;
assign feature_index_7[56] = 10'd101;
assign feature_index_7[57] = 10'd96;
assign feature_index_7[58] = 10'd270;
assign feature_index_7[59] = 10'd324;
assign feature_index_7[60] = 10'd216;
assign feature_index_7[61] = 10'd299;
assign feature_index_7[62] = 10'd564;
assign feature_index_7[63] = 10'd564;
assign feature_index_7[64] = 10'd265;
assign feature_index_7[65] = 10'd150;
assign feature_index_7[66] = 10'd358;
assign feature_index_7[67] = 10'd238;
assign feature_index_7[68] = 10'd376;
assign feature_index_7[69] = 10'd597;
assign feature_index_7[70] = 10'd0;
assign feature_index_7[71] = 10'd152;
assign feature_index_7[72] = 10'd513;
assign feature_index_7[73] = 10'd297;
assign feature_index_7[74] = 10'd513;
assign feature_index_7[75] = 10'd661;
assign feature_index_7[76] = 10'd376;
assign feature_index_7[77] = 10'd268;
assign feature_index_7[78] = 10'd485;
assign feature_index_7[79] = 10'd179;
assign feature_index_7[80] = 10'd382;
assign feature_index_7[81] = 10'd123;
assign feature_index_7[82] = 10'd385;
assign feature_index_7[83] = 10'd329;
assign feature_index_7[84] = 10'd625;
assign feature_index_7[85] = 10'd266;
assign feature_index_7[86] = 10'd329;
assign feature_index_7[87] = 10'd99;
assign feature_index_7[88] = 10'd563;
assign feature_index_7[89] = 10'd204;
assign feature_index_7[90] = 10'd239;
assign feature_index_7[91] = 10'd96;
assign feature_index_7[92] = 10'd628;
assign feature_index_7[93] = 10'd627;
assign feature_index_7[94] = 10'd454;
assign feature_index_7[95] = 10'd609;
assign feature_index_7[96] = 10'd407;
assign feature_index_7[97] = 10'd515;
assign feature_index_7[98] = 10'd658;
assign feature_index_7[99] = 10'd321;
assign feature_index_7[100] = 10'd372;
assign feature_index_7[101] = 10'd579;
assign feature_index_7[102] = 10'd262;
assign feature_index_7[103] = 10'd465;
assign feature_index_7[104] = 10'd566;
assign feature_index_7[105] = 10'd582;
assign feature_index_7[106] = 10'd316;
assign feature_index_7[107] = 10'd182;
assign feature_index_7[108] = 10'd315;
assign feature_index_7[109] = 10'd210;
assign feature_index_7[110] = 10'd683;
assign feature_index_7[111] = 10'd152;
assign feature_index_7[112] = 10'd545;
assign feature_index_7[113] = 10'd125;
assign feature_index_7[114] = 10'd188;
assign feature_index_7[115] = 10'd543;
assign feature_index_7[116] = 10'd577;
assign feature_index_7[117] = 10'd513;
assign feature_index_7[118] = 10'd318;
assign feature_index_7[119] = 10'd430;
assign feature_index_7[120] = 10'd294;
assign feature_index_7[121] = 10'd526;
assign feature_index_7[122] = 10'd0;
assign feature_index_7[123] = 10'd435;
assign feature_index_7[124] = 10'd245;
assign feature_index_7[125] = 10'd458;
assign feature_index_7[126] = 10'd573;
assign feature_index_7[127] = 10'd432;
assign feature_index_7[128] = 10'd215;
assign feature_index_7[129] = 10'd399;
assign feature_index_7[130] = 10'd378;
assign feature_index_7[131] = 10'd377;
assign feature_index_7[132] = 10'd210;
assign feature_index_7[133] = 10'd619;
assign feature_index_7[134] = 10'd205;
assign feature_index_7[135] = 10'd551;
assign feature_index_7[136] = 10'd132;
assign feature_index_7[137] = 10'd159;
assign feature_index_7[138] = 10'd401;
assign feature_index_7[139] = 10'd239;
assign feature_index_7[140] = 10'd429;
assign feature_index_7[141] = 10'd0;
assign feature_index_7[142] = 10'd0;
assign feature_index_7[143] = 10'd295;
assign feature_index_7[144] = 10'd487;
assign feature_index_7[145] = 10'd289;
assign feature_index_7[146] = 10'd153;
assign feature_index_7[147] = 10'd571;
assign feature_index_7[148] = 10'd485;
assign feature_index_7[149] = 10'd290;
assign feature_index_7[150] = 10'd603;
assign feature_index_7[151] = 10'd566;
assign feature_index_7[152] = 10'd497;
assign feature_index_7[153] = 10'd436;
assign feature_index_7[154] = 10'd458;
assign feature_index_7[155] = 10'd515;
assign feature_index_7[156] = 10'd656;
assign feature_index_7[157] = 10'd267;
assign feature_index_7[158] = 10'd659;
assign feature_index_7[159] = 10'd129;
assign feature_index_7[160] = 10'd512;
assign feature_index_7[161] = 10'd162;
assign feature_index_7[162] = 10'd325;
assign feature_index_7[163] = 10'd657;
assign feature_index_7[164] = 10'd321;
assign feature_index_7[165] = 10'd407;
assign feature_index_7[166] = 10'd149;
assign feature_index_7[167] = 10'd248;
assign feature_index_7[168] = 10'd354;
assign feature_index_7[169] = 10'd598;
assign feature_index_7[170] = 10'd462;
assign feature_index_7[171] = 10'd272;
assign feature_index_7[172] = 10'd124;
assign feature_index_7[173] = 10'd298;
assign feature_index_7[174] = 10'd547;
assign feature_index_7[175] = 10'd301;
assign feature_index_7[176] = 10'd242;
assign feature_index_7[177] = 10'd374;
assign feature_index_7[178] = 10'd0;
assign feature_index_7[179] = 10'd179;
assign feature_index_7[180] = 10'd492;
assign feature_index_7[181] = 10'd575;
assign feature_index_7[182] = 10'd292;
assign feature_index_7[183] = 10'd411;
assign feature_index_7[184] = 10'd397;
assign feature_index_7[185] = 10'd96;
assign feature_index_7[186] = 10'd145;
assign feature_index_7[187] = 10'd547;
assign feature_index_7[188] = 10'd271;
assign feature_index_7[189] = 10'd314;
assign feature_index_7[190] = 10'd265;
assign feature_index_7[191] = 10'd550;
assign feature_index_7[192] = 10'd466;
assign feature_index_7[193] = 10'd512;
assign feature_index_7[194] = 10'd122;
assign feature_index_7[195] = 10'd269;
assign feature_index_7[196] = 10'd569;
assign feature_index_7[197] = 10'd158;
assign feature_index_7[198] = 10'd325;
assign feature_index_7[199] = 10'd152;
assign feature_index_7[200] = 10'd267;
assign feature_index_7[201] = 10'd542;
assign feature_index_7[202] = 10'd498;
assign feature_index_7[203] = 10'd599;
assign feature_index_7[204] = 10'd330;
assign feature_index_7[205] = 10'd629;
assign feature_index_7[206] = 10'd464;
assign feature_index_7[207] = 10'd577;
assign feature_index_7[208] = 10'd265;
assign feature_index_7[209] = 10'd124;
assign feature_index_7[210] = 10'd543;
assign feature_index_7[211] = 10'd568;
assign feature_index_7[212] = 10'd681;
assign feature_index_7[213] = 10'd376;
assign feature_index_7[214] = 10'd153;
assign feature_index_7[215] = 10'd377;
assign feature_index_7[216] = 10'd371;
assign feature_index_7[217] = 10'd72;
assign feature_index_7[218] = 10'd213;
assign feature_index_7[219] = 10'd296;
assign feature_index_7[220] = 10'd466;
assign feature_index_7[221] = 10'd237;
assign feature_index_7[222] = 10'd229;
assign feature_index_7[223] = 10'd514;
assign feature_index_7[224] = 10'd379;
assign feature_index_7[225] = 10'd355;
assign feature_index_7[226] = 10'd214;
assign feature_index_7[227] = 10'd210;
assign feature_index_7[228] = 10'd545;
assign feature_index_7[229] = 10'd297;
assign feature_index_7[230] = 10'd550;
assign feature_index_7[231] = 10'd597;
assign feature_index_7[232] = 10'd429;
assign feature_index_7[233] = 10'd552;
assign feature_index_7[234] = 10'd213;
assign feature_index_7[235] = 10'd431;
assign feature_index_7[236] = 10'd639;
assign feature_index_7[237] = 10'd511;
assign feature_index_7[238] = 10'd499;
assign feature_index_7[239] = 10'd135;
assign feature_index_7[240] = 10'd0;
assign feature_index_7[241] = 10'd291;
assign feature_index_7[242] = 10'd493;
assign feature_index_7[243] = 10'd0;
assign feature_index_7[244] = 10'd441;
assign feature_index_7[245] = 10'd0;
assign feature_index_7[246] = 10'd0;
assign feature_index_7[247] = 10'd296;
assign feature_index_7[248] = 10'd468;
assign feature_index_7[249] = 10'd212;
assign feature_index_7[250] = 10'd0;
assign feature_index_7[251] = 10'd441;
assign feature_index_7[252] = 10'd74;
assign feature_index_7[253] = 10'd0;
assign feature_index_7[254] = 10'd403;
assign feature_index_7[255] = 10'd515;
assign feature_index_7[256] = 10'd626;
assign feature_index_7[257] = 10'd236;
assign feature_index_7[258] = 10'd396;
assign feature_index_7[259] = 10'd523;
assign feature_index_7[260] = 10'd327;
assign feature_index_7[261] = 10'd623;
assign feature_index_7[262] = 10'd321;
assign feature_index_7[263] = 10'd296;
assign feature_index_7[264] = 10'd240;
assign feature_index_7[265] = 10'd521;
assign feature_index_7[266] = 10'd239;
assign feature_index_7[267] = 10'd324;
assign feature_index_7[268] = 10'd408;
assign feature_index_7[269] = 10'd454;
assign feature_index_7[270] = 10'd563;
assign feature_index_7[271] = 10'd319;
assign feature_index_7[272] = 10'd245;
assign feature_index_7[273] = 10'd404;
assign feature_index_7[274] = 10'd353;
assign feature_index_7[275] = 10'd238;
assign feature_index_7[276] = 10'd570;
assign feature_index_7[277] = 10'd236;
assign feature_index_7[278] = 10'd327;
assign feature_index_7[279] = 10'd515;
assign feature_index_7[280] = 10'd551;
assign feature_index_7[281] = 10'd571;
assign feature_index_7[282] = 10'd404;
assign feature_index_7[283] = 10'd0;
assign feature_index_7[284] = 10'd0;
assign feature_index_7[285] = 10'd0;
assign feature_index_7[286] = 10'd0;
assign feature_index_7[287] = 10'd238;
assign feature_index_7[288] = 10'd376;
assign feature_index_7[289] = 10'd343;
assign feature_index_7[290] = 10'd98;
assign feature_index_7[291] = 10'd296;
assign feature_index_7[292] = 10'd346;
assign feature_index_7[293] = 10'd320;
assign feature_index_7[294] = 10'd298;
assign feature_index_7[295] = 10'd271;
assign feature_index_7[296] = 10'd299;
assign feature_index_7[297] = 10'd299;
assign feature_index_7[298] = 10'd264;
assign feature_index_7[299] = 10'd625;
assign feature_index_7[300] = 10'd653;
assign feature_index_7[301] = 10'd349;
assign feature_index_7[302] = 10'd318;
assign feature_index_7[303] = 10'd496;
assign feature_index_7[304] = 10'd487;
assign feature_index_7[305] = 10'd462;
assign feature_index_7[306] = 10'd351;
assign feature_index_7[307] = 10'd408;
assign feature_index_7[308] = 10'd324;
assign feature_index_7[309] = 10'd268;
assign feature_index_7[310] = 10'd241;
assign feature_index_7[311] = 10'd297;
assign feature_index_7[312] = 10'd182;
assign feature_index_7[313] = 10'd625;
assign feature_index_7[314] = 10'd487;
assign feature_index_7[315] = 10'd326;
assign feature_index_7[316] = 10'd628;
assign feature_index_7[317] = 10'd126;
assign feature_index_7[318] = 10'd270;
assign feature_index_7[319] = 10'd95;
assign feature_index_7[320] = 10'd375;
assign feature_index_7[321] = 10'd261;
assign feature_index_7[322] = 10'd350;
assign feature_index_7[323] = 10'd425;
assign feature_index_7[324] = 10'd326;
assign feature_index_7[325] = 10'd190;
assign feature_index_7[326] = 10'd487;
assign feature_index_7[327] = 10'd181;
assign feature_index_7[328] = 10'd457;
assign feature_index_7[329] = 10'd359;
assign feature_index_7[330] = 10'd431;
assign feature_index_7[331] = 10'd430;
assign feature_index_7[332] = 10'd318;
assign feature_index_7[333] = 10'd380;
assign feature_index_7[334] = 10'd628;
assign feature_index_7[335] = 10'd354;
assign feature_index_7[336] = 10'd360;
assign feature_index_7[337] = 10'd437;
assign feature_index_7[338] = 10'd0;
assign feature_index_7[339] = 10'd211;
assign feature_index_7[340] = 10'd462;
assign feature_index_7[341] = 10'd583;
assign feature_index_7[342] = 10'd434;
assign feature_index_7[343] = 10'd127;
assign feature_index_7[344] = 10'd354;
assign feature_index_7[345] = 10'd357;
assign feature_index_7[346] = 10'd295;
assign feature_index_7[347] = 10'd567;
assign feature_index_7[348] = 10'd275;
assign feature_index_7[349] = 10'd380;
assign feature_index_7[350] = 10'd152;
assign feature_index_7[351] = 10'd428;
assign feature_index_7[352] = 10'd488;
assign feature_index_7[353] = 10'd323;
assign feature_index_7[354] = 10'd462;
assign feature_index_7[355] = 10'd411;
assign feature_index_7[356] = 10'd406;
assign feature_index_7[357] = 10'd0;
assign feature_index_7[358] = 10'd0;
assign feature_index_7[359] = 10'd188;
assign feature_index_7[360] = 10'd654;
assign feature_index_7[361] = 10'd181;
assign feature_index_7[362] = 10'd471;
assign feature_index_7[363] = 10'd218;
assign feature_index_7[364] = 10'd455;
assign feature_index_7[365] = 10'd399;
assign feature_index_7[366] = 10'd563;
assign feature_index_7[367] = 10'd492;
assign feature_index_7[368] = 10'd185;
assign feature_index_7[369] = 10'd0;
assign feature_index_7[370] = 10'd0;
assign feature_index_7[371] = 10'd244;
assign feature_index_7[372] = 10'd0;
assign feature_index_7[373] = 10'd358;
assign feature_index_7[374] = 10'd330;
assign feature_index_7[375] = 10'd454;
assign feature_index_7[376] = 10'd135;
assign feature_index_7[377] = 10'd486;
assign feature_index_7[378] = 10'd237;
assign feature_index_7[379] = 10'd455;
assign feature_index_7[380] = 10'd403;
assign feature_index_7[381] = 10'd629;
assign feature_index_7[382] = 10'd174;
assign feature_index_7[383] = 10'd299;
assign feature_index_7[384] = 10'd487;
assign feature_index_7[385] = 10'd468;
assign feature_index_7[386] = 10'd428;
assign feature_index_7[387] = 10'd472;
assign feature_index_7[388] = 10'd242;
assign feature_index_7[389] = 10'd632;
assign feature_index_7[390] = 10'd540;
assign feature_index_7[391] = 10'd315;
assign feature_index_7[392] = 10'd655;
assign feature_index_7[393] = 10'd525;
assign feature_index_7[394] = 10'd155;
assign feature_index_7[395] = 10'd399;
assign feature_index_7[396] = 10'd494;
assign feature_index_7[397] = 10'd488;
assign feature_index_7[398] = 10'd440;
assign feature_index_7[399] = 10'd238;
assign feature_index_7[400] = 10'd543;
assign feature_index_7[401] = 10'd498;
assign feature_index_7[402] = 10'd260;
assign feature_index_7[403] = 10'd467;
assign feature_index_7[404] = 10'd320;
assign feature_index_7[405] = 10'd630;
assign feature_index_7[406] = 10'd603;
assign feature_index_7[407] = 10'd488;
assign feature_index_7[408] = 10'd688;
assign feature_index_7[409] = 10'd0;
assign feature_index_7[410] = 10'd0;
assign feature_index_7[411] = 10'd0;
assign feature_index_7[412] = 10'd708;
assign feature_index_7[413] = 10'd625;
assign feature_index_7[414] = 10'd661;
assign feature_index_7[415] = 10'd457;
assign feature_index_7[416] = 10'd543;
assign feature_index_7[417] = 10'd65;
assign feature_index_7[418] = 10'd399;
assign feature_index_7[419] = 10'd541;
assign feature_index_7[420] = 10'd262;
assign feature_index_7[421] = 10'd379;
assign feature_index_7[422] = 10'd0;
assign feature_index_7[423] = 10'd655;
assign feature_index_7[424] = 10'd349;
assign feature_index_7[425] = 10'd691;
assign feature_index_7[426] = 10'd230;
assign feature_index_7[427] = 10'd543;
assign feature_index_7[428] = 10'd556;
assign feature_index_7[429] = 10'd218;
assign feature_index_7[430] = 10'd99;
assign feature_index_7[431] = 10'd439;
assign feature_index_7[432] = 10'd457;
assign feature_index_7[433] = 10'd524;
assign feature_index_7[434] = 10'd354;
assign feature_index_7[435] = 10'd318;
assign feature_index_7[436] = 10'd441;
assign feature_index_7[437] = 10'd385;
assign feature_index_7[438] = 10'd660;
assign feature_index_7[439] = 10'd468;
assign feature_index_7[440] = 10'd290;
assign feature_index_7[441] = 10'd513;
assign feature_index_7[442] = 10'd625;
assign feature_index_7[443] = 10'd689;
assign feature_index_7[444] = 10'd178;
assign feature_index_7[445] = 10'd202;
assign feature_index_7[446] = 10'd467;
assign feature_index_7[447] = 10'd407;
assign feature_index_7[448] = 10'd429;
assign feature_index_7[449] = 10'd411;
assign feature_index_7[450] = 10'd467;
assign feature_index_7[451] = 10'd235;
assign feature_index_7[452] = 10'd100;
assign feature_index_7[453] = 10'd500;
assign feature_index_7[454] = 10'd551;
assign feature_index_7[455] = 10'd235;
assign feature_index_7[456] = 10'd213;
assign feature_index_7[457] = 10'd492;
assign feature_index_7[458] = 10'd243;
assign feature_index_7[459] = 10'd236;
assign feature_index_7[460] = 10'd626;
assign feature_index_7[461] = 10'd0;
assign feature_index_7[462] = 10'd452;
assign feature_index_7[463] = 10'd409;
assign feature_index_7[464] = 10'd486;
assign feature_index_7[465] = 10'd538;
assign feature_index_7[466] = 10'd658;
assign feature_index_7[467] = 10'd243;
assign feature_index_7[468] = 10'd120;
assign feature_index_7[469] = 10'd266;
assign feature_index_7[470] = 10'd627;
assign feature_index_7[471] = 10'd318;
assign feature_index_7[472] = 10'd398;
assign feature_index_7[473] = 10'd361;
assign feature_index_7[474] = 10'd0;
assign feature_index_7[475] = 10'd515;
assign feature_index_7[476] = 10'd0;
assign feature_index_7[477] = 10'd609;
assign feature_index_7[478] = 10'd567;
assign feature_index_7[479] = 10'd0;
assign feature_index_7[480] = 10'd0;
assign feature_index_7[481] = 10'd0;
assign feature_index_7[482] = 10'd0;
assign feature_index_7[483] = 10'd0;
assign feature_index_7[484] = 10'd0;
assign feature_index_7[485] = 10'd0;
assign feature_index_7[486] = 10'd0;
assign feature_index_7[487] = 10'd0;
assign feature_index_7[488] = 10'd0;
assign feature_index_7[489] = 10'd0;
assign feature_index_7[490] = 10'd0;
assign feature_index_7[491] = 10'd0;
assign feature_index_7[492] = 10'd0;
assign feature_index_7[493] = 10'd0;
assign feature_index_7[494] = 10'd0;
assign feature_index_7[495] = 10'd0;
assign feature_index_7[496] = 10'd0;
assign feature_index_7[497] = 10'd377;
assign feature_index_7[498] = 10'd0;
assign feature_index_7[499] = 10'd0;
assign feature_index_7[500] = 10'd0;
assign feature_index_7[501] = 10'd0;
assign feature_index_7[502] = 10'd0;
assign feature_index_7[503] = 10'd408;
assign feature_index_7[504] = 10'd0;
assign feature_index_7[505] = 10'd440;
assign feature_index_7[506] = 10'd0;
assign feature_index_7[507] = 10'd0;
assign feature_index_7[508] = 10'd0;
assign feature_index_7[509] = 10'd0;
assign feature_index_7[510] = 10'd272;
assign feature_index_7[511] = 10'd594;
assign feature_index_7[512] = 10'd385;
assign feature_index_7[513] = 10'd453;
assign feature_index_7[514] = 10'd243;
assign feature_index_7[515] = 10'd596;
assign feature_index_7[516] = 10'd0;
assign feature_index_7[517] = 10'd0;
assign feature_index_7[518] = 10'd291;
assign feature_index_7[519] = 10'd289;
assign feature_index_7[520] = 10'd479;
assign feature_index_7[521] = 10'd234;
assign feature_index_7[522] = 10'd237;
assign feature_index_7[523] = 10'd459;
assign feature_index_7[524] = 10'd149;
assign feature_index_7[525] = 10'd523;
assign feature_index_7[526] = 10'd380;
assign feature_index_7[527] = 10'd596;
assign feature_index_7[528] = 10'd291;
assign feature_index_7[529] = 10'd184;
assign feature_index_7[530] = 10'd518;
assign feature_index_7[531] = 10'd489;
assign feature_index_7[532] = 10'd378;
assign feature_index_7[533] = 10'd298;
assign feature_index_7[534] = 10'd202;
assign feature_index_7[535] = 10'd179;
assign feature_index_7[536] = 10'd320;
assign feature_index_7[537] = 10'd161;
assign feature_index_7[538] = 10'd343;
assign feature_index_7[539] = 10'd577;
assign feature_index_7[540] = 10'd510;
assign feature_index_7[541] = 10'd0;
assign feature_index_7[542] = 10'd0;
assign feature_index_7[543] = 10'd298;
assign feature_index_7[544] = 10'd495;
assign feature_index_7[545] = 10'd469;
assign feature_index_7[546] = 10'd599;
assign feature_index_7[547] = 10'd571;
assign feature_index_7[548] = 10'd236;
assign feature_index_7[549] = 10'd268;
assign feature_index_7[550] = 10'd571;
assign feature_index_7[551] = 10'd210;
assign feature_index_7[552] = 10'd153;
assign feature_index_7[553] = 10'd464;
assign feature_index_7[554] = 10'd490;
assign feature_index_7[555] = 10'd684;
assign feature_index_7[556] = 10'd483;
assign feature_index_7[557] = 10'd202;
assign feature_index_7[558] = 10'd601;
assign feature_index_7[559] = 10'd241;
assign feature_index_7[560] = 10'd634;
assign feature_index_7[561] = 10'd0;
assign feature_index_7[562] = 10'd122;
assign feature_index_7[563] = 10'd0;
assign feature_index_7[564] = 10'd0;
assign feature_index_7[565] = 10'd408;
assign feature_index_7[566] = 10'd0;
assign feature_index_7[567] = 10'd0;
assign feature_index_7[568] = 10'd0;
assign feature_index_7[569] = 10'd0;
assign feature_index_7[570] = 10'd0;
assign feature_index_7[571] = 10'd0;
assign feature_index_7[572] = 10'd0;
assign feature_index_7[573] = 10'd0;
assign feature_index_7[574] = 10'd0;
assign feature_index_7[575] = 10'd536;
assign feature_index_7[576] = 10'd567;
assign feature_index_7[577] = 10'd490;
assign feature_index_7[578] = 10'd289;
assign feature_index_7[579] = 10'd518;
assign feature_index_7[580] = 10'd242;
assign feature_index_7[581] = 10'd659;
assign feature_index_7[582] = 10'd208;
assign feature_index_7[583] = 10'd518;
assign feature_index_7[584] = 10'd375;
assign feature_index_7[585] = 10'd299;
assign feature_index_7[586] = 10'd265;
assign feature_index_7[587] = 10'd0;
assign feature_index_7[588] = 10'd218;
assign feature_index_7[589] = 10'd287;
assign feature_index_7[590] = 10'd347;
assign feature_index_7[591] = 10'd543;
assign feature_index_7[592] = 10'd412;
assign feature_index_7[593] = 10'd659;
assign feature_index_7[594] = 10'd378;
assign feature_index_7[595] = 10'd435;
assign feature_index_7[596] = 10'd351;
assign feature_index_7[597] = 10'd554;
assign feature_index_7[598] = 10'd569;
assign feature_index_7[599] = 10'd439;
assign feature_index_7[600] = 10'd348;
assign feature_index_7[601] = 10'd266;
assign feature_index_7[602] = 10'd161;
assign feature_index_7[603] = 10'd685;
assign feature_index_7[604] = 10'd0;
assign feature_index_7[605] = 10'd350;
assign feature_index_7[606] = 10'd352;
assign feature_index_7[607] = 10'd609;
assign feature_index_7[608] = 10'd244;
assign feature_index_7[609] = 10'd0;
assign feature_index_7[610] = 10'd0;
assign feature_index_7[611] = 10'd493;
assign feature_index_7[612] = 10'd660;
assign feature_index_7[613] = 10'd271;
assign feature_index_7[614] = 10'd209;
assign feature_index_7[615] = 10'd349;
assign feature_index_7[616] = 10'd0;
assign feature_index_7[617] = 10'd435;
assign feature_index_7[618] = 10'd517;
assign feature_index_7[619] = 10'd185;
assign feature_index_7[620] = 10'd295;
assign feature_index_7[621] = 10'd100;
assign feature_index_7[622] = 10'd570;
assign feature_index_7[623] = 10'd632;
assign feature_index_7[624] = 10'd653;
assign feature_index_7[625] = 10'd459;
assign feature_index_7[626] = 10'd214;
assign feature_index_7[627] = 10'd484;
assign feature_index_7[628] = 10'd151;
assign feature_index_7[629] = 10'd154;
assign feature_index_7[630] = 10'd262;
assign feature_index_7[631] = 10'd519;
assign feature_index_7[632] = 10'd413;
assign feature_index_7[633] = 10'd666;
assign feature_index_7[634] = 10'd564;
assign feature_index_7[635] = 10'd443;
assign feature_index_7[636] = 10'd239;
assign feature_index_7[637] = 10'd491;
assign feature_index_7[638] = 10'd329;
assign feature_index_7[639] = 10'd479;
assign feature_index_7[640] = 10'd294;
assign feature_index_7[641] = 10'd513;
assign feature_index_7[642] = 10'd126;
assign feature_index_7[643] = 10'd490;
assign feature_index_7[644] = 10'd514;
assign feature_index_7[645] = 10'd157;
assign feature_index_7[646] = 10'd207;
assign feature_index_7[647] = 10'd263;
assign feature_index_7[648] = 10'd540;
assign feature_index_7[649] = 10'd313;
assign feature_index_7[650] = 10'd380;
assign feature_index_7[651] = 10'd235;
assign feature_index_7[652] = 10'd229;
assign feature_index_7[653] = 10'd164;
assign feature_index_7[654] = 10'd517;
assign feature_index_7[655] = 10'd352;
assign feature_index_7[656] = 10'd325;
assign feature_index_7[657] = 10'd545;
assign feature_index_7[658] = 10'd325;
assign feature_index_7[659] = 10'd432;
assign feature_index_7[660] = 10'd0;
assign feature_index_7[661] = 10'd262;
assign feature_index_7[662] = 10'd435;
assign feature_index_7[663] = 10'd657;
assign feature_index_7[664] = 10'd327;
assign feature_index_7[665] = 10'd177;
assign feature_index_7[666] = 10'd298;
assign feature_index_7[667] = 10'd102;
assign feature_index_7[668] = 10'd180;
assign feature_index_7[669] = 10'd0;
assign feature_index_7[670] = 10'd0;
assign feature_index_7[671] = 10'd582;
assign feature_index_7[672] = 10'd290;
assign feature_index_7[673] = 10'd526;
assign feature_index_7[674] = 10'd0;
assign feature_index_7[675] = 10'd0;
assign feature_index_7[676] = 10'd295;
assign feature_index_7[677] = 10'd0;
assign feature_index_7[678] = 10'd0;
assign feature_index_7[679] = 10'd512;
assign feature_index_7[680] = 10'd566;
assign feature_index_7[681] = 10'd627;
assign feature_index_7[682] = 10'd541;
assign feature_index_7[683] = 10'd553;
assign feature_index_7[684] = 10'd0;
assign feature_index_7[685] = 10'd0;
assign feature_index_7[686] = 10'd492;
assign feature_index_7[687] = 10'd291;
assign feature_index_7[688] = 10'd268;
assign feature_index_7[689] = 10'd276;
assign feature_index_7[690] = 10'd455;
assign feature_index_7[691] = 10'd175;
assign feature_index_7[692] = 10'd206;
assign feature_index_7[693] = 10'd509;
assign feature_index_7[694] = 10'd231;
assign feature_index_7[695] = 10'd570;
assign feature_index_7[696] = 10'd626;
assign feature_index_7[697] = 10'd512;
assign feature_index_7[698] = 10'd0;
assign feature_index_7[699] = 10'd149;
assign feature_index_7[700] = 10'd595;
assign feature_index_7[701] = 10'd384;
assign feature_index_7[702] = 10'd240;
assign feature_index_7[703] = 10'd565;
assign feature_index_7[704] = 10'd103;
assign feature_index_7[705] = 10'd201;
assign feature_index_7[706] = 10'd149;
assign feature_index_7[707] = 10'd69;
assign feature_index_7[708] = 10'd326;
assign feature_index_7[709] = 10'd0;
assign feature_index_7[710] = 10'd0;
assign feature_index_7[711] = 10'd93;
assign feature_index_7[712] = 10'd654;
assign feature_index_7[713] = 10'd0;
assign feature_index_7[714] = 10'd574;
assign feature_index_7[715] = 10'd0;
assign feature_index_7[716] = 10'd0;
assign feature_index_7[717] = 10'd0;
assign feature_index_7[718] = 10'd0;
assign feature_index_7[719] = 10'd128;
assign feature_index_7[720] = 10'd270;
assign feature_index_7[721] = 10'd553;
assign feature_index_7[722] = 10'd317;
assign feature_index_7[723] = 10'd122;
assign feature_index_7[724] = 10'd214;
assign feature_index_7[725] = 10'd487;
assign feature_index_7[726] = 10'd0;
assign feature_index_7[727] = 10'd554;
assign feature_index_7[728] = 10'd581;
assign feature_index_7[729] = 10'd0;
assign feature_index_7[730] = 10'd627;
assign feature_index_7[731] = 10'd381;
assign feature_index_7[732] = 10'd609;
assign feature_index_7[733] = 10'd408;
assign feature_index_7[734] = 10'd0;
assign feature_index_7[735] = 10'd576;
assign feature_index_7[736] = 10'd609;
assign feature_index_7[737] = 10'd286;
assign feature_index_7[738] = 10'd593;
assign feature_index_7[739] = 10'd0;
assign feature_index_7[740] = 10'd0;
assign feature_index_7[741] = 10'd0;
assign feature_index_7[742] = 10'd0;
assign feature_index_7[743] = 10'd266;
assign feature_index_7[744] = 10'd638;
assign feature_index_7[745] = 10'd0;
assign feature_index_7[746] = 10'd0;
assign feature_index_7[747] = 10'd102;
assign feature_index_7[748] = 10'd216;
assign feature_index_7[749] = 10'd189;
assign feature_index_7[750] = 10'd552;
assign feature_index_7[751] = 10'd0;
assign feature_index_7[752] = 10'd0;
assign feature_index_7[753] = 10'd0;
assign feature_index_7[754] = 10'd0;
assign feature_index_7[755] = 10'd574;
assign feature_index_7[756] = 10'd500;
assign feature_index_7[757] = 10'd522;
assign feature_index_7[758] = 10'd275;
assign feature_index_7[759] = 10'd270;
assign feature_index_7[760] = 10'd267;
assign feature_index_7[761] = 10'd416;
assign feature_index_7[762] = 10'd348;
assign feature_index_7[763] = 10'd404;
assign feature_index_7[764] = 10'd184;
assign feature_index_7[765] = 10'd131;
assign feature_index_7[766] = 10'd663;
assign feature_index_7[767] = 10'd206;
assign feature_index_7[768] = 10'd602;
assign feature_index_7[769] = 10'd399;
assign feature_index_7[770] = 10'd321;
assign feature_index_7[771] = 10'd385;
assign feature_index_7[772] = 10'd0;
assign feature_index_7[773] = 10'd0;
assign feature_index_7[774] = 10'd0;
assign feature_index_7[775] = 10'd664;
assign feature_index_7[776] = 10'd0;
assign feature_index_7[777] = 10'd570;
assign feature_index_7[778] = 10'd636;
assign feature_index_7[779] = 10'd576;
assign feature_index_7[780] = 10'd375;
assign feature_index_7[781] = 10'd0;
assign feature_index_7[782] = 10'd0;
assign feature_index_7[783] = 10'd518;
assign feature_index_7[784] = 10'd353;
assign feature_index_7[785] = 10'd386;
assign feature_index_7[786] = 10'd516;
assign feature_index_7[787] = 10'd659;
assign feature_index_7[788] = 10'd455;
assign feature_index_7[789] = 10'd238;
assign feature_index_7[790] = 10'd632;
assign feature_index_7[791] = 10'd441;
assign feature_index_7[792] = 10'd345;
assign feature_index_7[793] = 10'd206;
assign feature_index_7[794] = 10'd385;
assign feature_index_7[795] = 10'd320;
assign feature_index_7[796] = 10'd217;
assign feature_index_7[797] = 10'd317;
assign feature_index_7[798] = 10'd268;
assign feature_index_7[799] = 10'd465;
assign feature_index_7[800] = 10'd317;
assign feature_index_7[801] = 10'd210;
assign feature_index_7[802] = 10'd415;
assign feature_index_7[803] = 10'd407;
assign feature_index_7[804] = 10'd288;
assign feature_index_7[805] = 10'd382;
assign feature_index_7[806] = 10'd296;
assign feature_index_7[807] = 10'd688;
assign feature_index_7[808] = 10'd434;
assign feature_index_7[809] = 10'd370;
assign feature_index_7[810] = 10'd433;
assign feature_index_7[811] = 10'd654;
assign feature_index_7[812] = 10'd540;
assign feature_index_7[813] = 10'd238;
assign feature_index_7[814] = 10'd376;
assign feature_index_7[815] = 10'd593;
assign feature_index_7[816] = 10'd514;
assign feature_index_7[817] = 10'd262;
assign feature_index_7[818] = 10'd629;
assign feature_index_7[819] = 10'd0;
assign feature_index_7[820] = 10'd0;
assign feature_index_7[821] = 10'd0;
assign feature_index_7[822] = 10'd0;
assign feature_index_7[823] = 10'd0;
assign feature_index_7[824] = 10'd0;
assign feature_index_7[825] = 10'd0;
assign feature_index_7[826] = 10'd0;
assign feature_index_7[827] = 10'd0;
assign feature_index_7[828] = 10'd441;
assign feature_index_7[829] = 10'd573;
assign feature_index_7[830] = 10'd272;
assign feature_index_7[831] = 10'd653;
assign feature_index_7[832] = 10'd409;
assign feature_index_7[833] = 10'd328;
assign feature_index_7[834] = 10'd565;
assign feature_index_7[835] = 10'd94;
assign feature_index_7[836] = 10'd0;
assign feature_index_7[837] = 10'd260;
assign feature_index_7[838] = 10'd692;
assign feature_index_7[839] = 10'd371;
assign feature_index_7[840] = 10'd626;
assign feature_index_7[841] = 10'd385;
assign feature_index_7[842] = 10'd525;
assign feature_index_7[843] = 10'd257;
assign feature_index_7[844] = 10'd409;
assign feature_index_7[845] = 10'd0;
assign feature_index_7[846] = 10'd0;
assign feature_index_7[847] = 10'd376;
assign feature_index_7[848] = 10'd577;
assign feature_index_7[849] = 10'd595;
assign feature_index_7[850] = 10'd542;
assign feature_index_7[851] = 10'd314;
assign feature_index_7[852] = 10'd144;
assign feature_index_7[853] = 10'd668;
assign feature_index_7[854] = 10'd0;
assign feature_index_7[855] = 10'd373;
assign feature_index_7[856] = 10'd553;
assign feature_index_7[857] = 10'd346;
assign feature_index_7[858] = 10'd0;
assign feature_index_7[859] = 10'd410;
assign feature_index_7[860] = 10'd437;
assign feature_index_7[861] = 10'd456;
assign feature_index_7[862] = 10'd351;
assign feature_index_7[863] = 10'd220;
assign feature_index_7[864] = 10'd398;
assign feature_index_7[865] = 10'd521;
assign feature_index_7[866] = 10'd547;
assign feature_index_7[867] = 10'd379;
assign feature_index_7[868] = 10'd546;
assign feature_index_7[869] = 10'd433;
assign feature_index_7[870] = 10'd455;
assign feature_index_7[871] = 10'd192;
assign feature_index_7[872] = 10'd102;
assign feature_index_7[873] = 10'd345;
assign feature_index_7[874] = 10'd316;
assign feature_index_7[875] = 10'd514;
assign feature_index_7[876] = 10'd0;
assign feature_index_7[877] = 10'd469;
assign feature_index_7[878] = 10'd574;
assign feature_index_7[879] = 10'd494;
assign feature_index_7[880] = 10'd208;
assign feature_index_7[881] = 10'd246;
assign feature_index_7[882] = 10'd495;
assign feature_index_7[883] = 10'd331;
assign feature_index_7[884] = 10'd495;
assign feature_index_7[885] = 10'd579;
assign feature_index_7[886] = 10'd193;
assign feature_index_7[887] = 10'd346;
assign feature_index_7[888] = 10'd0;
assign feature_index_7[889] = 10'd352;
assign feature_index_7[890] = 10'd400;
assign feature_index_7[891] = 10'd481;
assign feature_index_7[892] = 10'd655;
assign feature_index_7[893] = 10'd0;
assign feature_index_7[894] = 10'd526;
assign feature_index_7[895] = 10'd408;
assign feature_index_7[896] = 10'd183;
assign feature_index_7[897] = 10'd128;
assign feature_index_7[898] = 10'd381;
assign feature_index_7[899] = 10'd322;
assign feature_index_7[900] = 10'd0;
assign feature_index_7[901] = 10'd491;
assign feature_index_7[902] = 10'd0;
assign feature_index_7[903] = 10'd516;
assign feature_index_7[904] = 10'd443;
assign feature_index_7[905] = 10'd326;
assign feature_index_7[906] = 10'd0;
assign feature_index_7[907] = 10'd527;
assign feature_index_7[908] = 10'd0;
assign feature_index_7[909] = 10'd629;
assign feature_index_7[910] = 10'd402;
assign feature_index_7[911] = 10'd680;
assign feature_index_7[912] = 10'd737;
assign feature_index_7[913] = 10'd428;
assign feature_index_7[914] = 10'd382;
assign feature_index_7[915] = 10'd547;
assign feature_index_7[916] = 10'd628;
assign feature_index_7[917] = 10'd657;
assign feature_index_7[918] = 10'd458;
assign feature_index_7[919] = 10'd571;
assign feature_index_7[920] = 10'd0;
assign feature_index_7[921] = 10'd0;
assign feature_index_7[922] = 10'd0;
assign feature_index_7[923] = 10'd0;
assign feature_index_7[924] = 10'd0;
assign feature_index_7[925] = 10'd0;
assign feature_index_7[926] = 10'd0;
assign feature_index_7[927] = 10'd655;
assign feature_index_7[928] = 10'd154;
assign feature_index_7[929] = 10'd352;
assign feature_index_7[930] = 10'd301;
assign feature_index_7[931] = 10'd514;
assign feature_index_7[932] = 10'd357;
assign feature_index_7[933] = 10'd99;
assign feature_index_7[934] = 10'd514;
assign feature_index_7[935] = 10'd0;
assign feature_index_7[936] = 10'd0;
assign feature_index_7[937] = 10'd0;
assign feature_index_7[938] = 10'd0;
assign feature_index_7[939] = 10'd230;
assign feature_index_7[940] = 10'd467;
assign feature_index_7[941] = 10'd0;
assign feature_index_7[942] = 10'd607;
assign feature_index_7[943] = 10'd524;
assign feature_index_7[944] = 10'd403;
assign feature_index_7[945] = 10'd268;
assign feature_index_7[946] = 10'd380;
assign feature_index_7[947] = 10'd149;
assign feature_index_7[948] = 10'd0;
assign feature_index_7[949] = 10'd0;
assign feature_index_7[950] = 10'd0;
assign feature_index_7[951] = 10'd0;
assign feature_index_7[952] = 10'd156;
assign feature_index_7[953] = 10'd0;
assign feature_index_7[954] = 10'd0;
assign feature_index_7[955] = 10'd379;
assign feature_index_7[956] = 10'd0;
assign feature_index_7[957] = 10'd0;
assign feature_index_7[958] = 10'd0;
assign feature_index_7[959] = 10'd0;
assign feature_index_7[960] = 10'd0;
assign feature_index_7[961] = 10'd0;
assign feature_index_7[962] = 10'd0;
assign feature_index_7[963] = 10'd0;
assign feature_index_7[964] = 10'd0;
assign feature_index_7[965] = 10'd0;
assign feature_index_7[966] = 10'd0;
assign feature_index_7[967] = 10'd0;
assign feature_index_7[968] = 10'd0;
assign feature_index_7[969] = 10'd0;
assign feature_index_7[970] = 10'd0;
assign feature_index_7[971] = 10'd0;
assign feature_index_7[972] = 10'd0;
assign feature_index_7[973] = 10'd0;
assign feature_index_7[974] = 10'd0;
assign feature_index_7[975] = 10'd0;
assign feature_index_7[976] = 10'd0;
assign feature_index_7[977] = 10'd0;
assign feature_index_7[978] = 10'd0;
assign feature_index_7[979] = 10'd0;
assign feature_index_7[980] = 10'd0;
assign feature_index_7[981] = 10'd0;
assign feature_index_7[982] = 10'd0;
assign feature_index_7[983] = 10'd0;
assign feature_index_7[984] = 10'd0;
assign feature_index_7[985] = 10'd0;
assign feature_index_7[986] = 10'd0;
assign feature_index_7[987] = 10'd0;
assign feature_index_7[988] = 10'd0;
assign feature_index_7[989] = 10'd0;
assign feature_index_7[990] = 10'd0;
assign feature_index_7[991] = 10'd0;
assign feature_index_7[992] = 10'd0;
assign feature_index_7[993] = 10'd0;
assign feature_index_7[994] = 10'd0;
assign feature_index_7[995] = 10'd0;
assign feature_index_7[996] = 10'd487;
assign feature_index_7[997] = 10'd0;
assign feature_index_7[998] = 10'd0;
assign feature_index_7[999] = 10'd0;
assign feature_index_7[1000] = 10'd0;
assign feature_index_7[1001] = 10'd0;
assign feature_index_7[1002] = 10'd0;
assign feature_index_7[1003] = 10'd0;
assign feature_index_7[1004] = 10'd0;
assign feature_index_7[1005] = 10'd0;
assign feature_index_7[1006] = 10'd0;
assign feature_index_7[1007] = 10'd0;
assign feature_index_7[1008] = 10'd574;
assign feature_index_7[1009] = 10'd0;
assign feature_index_7[1010] = 10'd0;
assign feature_index_7[1011] = 10'd566;
assign feature_index_7[1012] = 10'd0;
assign feature_index_7[1013] = 10'd0;
assign feature_index_7[1014] = 10'd0;
assign feature_index_7[1015] = 10'd0;
assign feature_index_7[1016] = 10'd0;
assign feature_index_7[1017] = 10'd0;
assign feature_index_7[1018] = 10'd0;
assign feature_index_7[1019] = 10'd0;
assign feature_index_7[1020] = 10'd0;
assign feature_index_7[1021] = 10'd0;
assign feature_index_7[1022] = 10'd0;
assign feature_index_8[0] = 10'd456;
assign feature_index_8[1] = 10'd346;
assign feature_index_8[2] = 10'd543;
assign feature_index_8[3] = 10'd550;
assign feature_index_8[4] = 10'd459;
assign feature_index_8[5] = 10'd628;
assign feature_index_8[6] = 10'd270;
assign feature_index_8[7] = 10'd264;
assign feature_index_8[8] = 10'd461;
assign feature_index_8[9] = 10'd468;
assign feature_index_8[10] = 10'd514;
assign feature_index_8[11] = 10'd182;
assign feature_index_8[12] = 10'd405;
assign feature_index_8[13] = 10'd215;
assign feature_index_8[14] = 10'd463;
assign feature_index_8[15] = 10'd351;
assign feature_index_8[16] = 10'd182;
assign feature_index_8[17] = 10'd343;
assign feature_index_8[18] = 10'd569;
assign feature_index_8[19] = 10'd184;
assign feature_index_8[20] = 10'd149;
assign feature_index_8[21] = 10'd653;
assign feature_index_8[22] = 10'd430;
assign feature_index_8[23] = 10'd149;
assign feature_index_8[24] = 10'd683;
assign feature_index_8[25] = 10'd464;
assign feature_index_8[26] = 10'd127;
assign feature_index_8[27] = 10'd602;
assign feature_index_8[28] = 10'd347;
assign feature_index_8[29] = 10'd373;
assign feature_index_8[30] = 10'd569;
assign feature_index_8[31] = 10'd154;
assign feature_index_8[32] = 10'd402;
assign feature_index_8[33] = 10'd381;
assign feature_index_8[34] = 10'd625;
assign feature_index_8[35] = 10'd627;
assign feature_index_8[36] = 10'd387;
assign feature_index_8[37] = 10'd681;
assign feature_index_8[38] = 10'd657;
assign feature_index_8[39] = 10'd567;
assign feature_index_8[40] = 10'd568;
assign feature_index_8[41] = 10'd350;
assign feature_index_8[42] = 10'd260;
assign feature_index_8[43] = 10'd239;
assign feature_index_8[44] = 10'd300;
assign feature_index_8[45] = 10'd293;
assign feature_index_8[46] = 10'd300;
assign feature_index_8[47] = 10'd186;
assign feature_index_8[48] = 10'd344;
assign feature_index_8[49] = 10'd289;
assign feature_index_8[50] = 10'd432;
assign feature_index_8[51] = 10'd461;
assign feature_index_8[52] = 10'd186;
assign feature_index_8[53] = 10'd317;
assign feature_index_8[54] = 10'd522;
assign feature_index_8[55] = 10'd574;
assign feature_index_8[56] = 10'd247;
assign feature_index_8[57] = 10'd315;
assign feature_index_8[58] = 10'd245;
assign feature_index_8[59] = 10'd399;
assign feature_index_8[60] = 10'd405;
assign feature_index_8[61] = 10'd211;
assign feature_index_8[62] = 10'd374;
assign feature_index_8[63] = 10'd158;
assign feature_index_8[64] = 10'd454;
assign feature_index_8[65] = 10'd465;
assign feature_index_8[66] = 10'd486;
assign feature_index_8[67] = 10'd349;
assign feature_index_8[68] = 10'd432;
assign feature_index_8[69] = 10'd214;
assign feature_index_8[70] = 10'd157;
assign feature_index_8[71] = 10'd262;
assign feature_index_8[72] = 10'd322;
assign feature_index_8[73] = 10'd434;
assign feature_index_8[74] = 10'd567;
assign feature_index_8[75] = 10'd544;
assign feature_index_8[76] = 10'd183;
assign feature_index_8[77] = 10'd319;
assign feature_index_8[78] = 10'd293;
assign feature_index_8[79] = 10'd321;
assign feature_index_8[80] = 10'd247;
assign feature_index_8[81] = 10'd155;
assign feature_index_8[82] = 10'd297;
assign feature_index_8[83] = 10'd510;
assign feature_index_8[84] = 10'd297;
assign feature_index_8[85] = 10'd368;
assign feature_index_8[86] = 10'd342;
assign feature_index_8[87] = 10'd543;
assign feature_index_8[88] = 10'd156;
assign feature_index_8[89] = 10'd153;
assign feature_index_8[90] = 10'd381;
assign feature_index_8[91] = 10'd683;
assign feature_index_8[92] = 10'd552;
assign feature_index_8[93] = 10'd99;
assign feature_index_8[94] = 10'd214;
assign feature_index_8[95] = 10'd269;
assign feature_index_8[96] = 10'd626;
assign feature_index_8[97] = 10'd569;
assign feature_index_8[98] = 10'd545;
assign feature_index_8[99] = 10'd347;
assign feature_index_8[100] = 10'd443;
assign feature_index_8[101] = 10'd350;
assign feature_index_8[102] = 10'd264;
assign feature_index_8[103] = 10'd353;
assign feature_index_8[104] = 10'd345;
assign feature_index_8[105] = 10'd460;
assign feature_index_8[106] = 10'd319;
assign feature_index_8[107] = 10'd180;
assign feature_index_8[108] = 10'd546;
assign feature_index_8[109] = 10'd373;
assign feature_index_8[110] = 10'd658;
assign feature_index_8[111] = 10'd681;
assign feature_index_8[112] = 10'd520;
assign feature_index_8[113] = 10'd621;
assign feature_index_8[114] = 10'd415;
assign feature_index_8[115] = 10'd319;
assign feature_index_8[116] = 10'd387;
assign feature_index_8[117] = 10'd232;
assign feature_index_8[118] = 10'd329;
assign feature_index_8[119] = 10'd431;
assign feature_index_8[120] = 10'd350;
assign feature_index_8[121] = 10'd440;
assign feature_index_8[122] = 10'd241;
assign feature_index_8[123] = 10'd353;
assign feature_index_8[124] = 10'd156;
assign feature_index_8[125] = 10'd349;
assign feature_index_8[126] = 10'd320;
assign feature_index_8[127] = 10'd241;
assign feature_index_8[128] = 10'd215;
assign feature_index_8[129] = 10'd635;
assign feature_index_8[130] = 10'd435;
assign feature_index_8[131] = 10'd178;
assign feature_index_8[132] = 10'd488;
assign feature_index_8[133] = 10'd344;
assign feature_index_8[134] = 10'd153;
assign feature_index_8[135] = 10'd401;
assign feature_index_8[136] = 10'd623;
assign feature_index_8[137] = 10'd125;
assign feature_index_8[138] = 10'd595;
assign feature_index_8[139] = 10'd234;
assign feature_index_8[140] = 10'd405;
assign feature_index_8[141] = 10'd482;
assign feature_index_8[142] = 10'd377;
assign feature_index_8[143] = 10'd178;
assign feature_index_8[144] = 10'd285;
assign feature_index_8[145] = 10'd378;
assign feature_index_8[146] = 10'd459;
assign feature_index_8[147] = 10'd655;
assign feature_index_8[148] = 10'd247;
assign feature_index_8[149] = 10'd208;
assign feature_index_8[150] = 10'd566;
assign feature_index_8[151] = 10'd429;
assign feature_index_8[152] = 10'd375;
assign feature_index_8[153] = 10'd409;
assign feature_index_8[154] = 10'd189;
assign feature_index_8[155] = 10'd357;
assign feature_index_8[156] = 10'd440;
assign feature_index_8[157] = 10'd124;
assign feature_index_8[158] = 10'd374;
assign feature_index_8[159] = 10'd209;
assign feature_index_8[160] = 10'd382;
assign feature_index_8[161] = 10'd414;
assign feature_index_8[162] = 10'd426;
assign feature_index_8[163] = 10'd546;
assign feature_index_8[164] = 10'd565;
assign feature_index_8[165] = 10'd331;
assign feature_index_8[166] = 10'd292;
assign feature_index_8[167] = 10'd374;
assign feature_index_8[168] = 10'd576;
assign feature_index_8[169] = 10'd328;
assign feature_index_8[170] = 10'd623;
assign feature_index_8[171] = 10'd146;
assign feature_index_8[172] = 10'd340;
assign feature_index_8[173] = 10'd267;
assign feature_index_8[174] = 10'd654;
assign feature_index_8[175] = 10'd237;
assign feature_index_8[176] = 10'd242;
assign feature_index_8[177] = 10'd626;
assign feature_index_8[178] = 10'd182;
assign feature_index_8[179] = 10'd516;
assign feature_index_8[180] = 10'd177;
assign feature_index_8[181] = 10'd152;
assign feature_index_8[182] = 10'd577;
assign feature_index_8[183] = 10'd348;
assign feature_index_8[184] = 10'd375;
assign feature_index_8[185] = 10'd658;
assign feature_index_8[186] = 10'd524;
assign feature_index_8[187] = 10'd544;
assign feature_index_8[188] = 10'd298;
assign feature_index_8[189] = 10'd183;
assign feature_index_8[190] = 10'd494;
assign feature_index_8[191] = 10'd238;
assign feature_index_8[192] = 10'd436;
assign feature_index_8[193] = 10'd274;
assign feature_index_8[194] = 10'd329;
assign feature_index_8[195] = 10'd210;
assign feature_index_8[196] = 10'd0;
assign feature_index_8[197] = 10'd296;
assign feature_index_8[198] = 10'd493;
assign feature_index_8[199] = 10'd286;
assign feature_index_8[200] = 10'd572;
assign feature_index_8[201] = 10'd382;
assign feature_index_8[202] = 10'd493;
assign feature_index_8[203] = 10'd437;
assign feature_index_8[204] = 10'd268;
assign feature_index_8[205] = 10'd155;
assign feature_index_8[206] = 10'd510;
assign feature_index_8[207] = 10'd518;
assign feature_index_8[208] = 10'd322;
assign feature_index_8[209] = 10'd383;
assign feature_index_8[210] = 10'd484;
assign feature_index_8[211] = 10'd569;
assign feature_index_8[212] = 10'd597;
assign feature_index_8[213] = 10'd521;
assign feature_index_8[214] = 10'd625;
assign feature_index_8[215] = 10'd212;
assign feature_index_8[216] = 10'd247;
assign feature_index_8[217] = 10'd511;
assign feature_index_8[218] = 10'd190;
assign feature_index_8[219] = 10'd439;
assign feature_index_8[220] = 10'd548;
assign feature_index_8[221] = 10'd291;
assign feature_index_8[222] = 10'd264;
assign feature_index_8[223] = 10'd327;
assign feature_index_8[224] = 10'd273;
assign feature_index_8[225] = 10'd273;
assign feature_index_8[226] = 10'd245;
assign feature_index_8[227] = 10'd685;
assign feature_index_8[228] = 10'd0;
assign feature_index_8[229] = 10'd410;
assign feature_index_8[230] = 10'd405;
assign feature_index_8[231] = 10'd349;
assign feature_index_8[232] = 10'd126;
assign feature_index_8[233] = 10'd511;
assign feature_index_8[234] = 10'd463;
assign feature_index_8[235] = 10'd485;
assign feature_index_8[236] = 10'd569;
assign feature_index_8[237] = 10'd387;
assign feature_index_8[238] = 10'd353;
assign feature_index_8[239] = 10'd595;
assign feature_index_8[240] = 10'd346;
assign feature_index_8[241] = 10'd629;
assign feature_index_8[242] = 10'd120;
assign feature_index_8[243] = 10'd442;
assign feature_index_8[244] = 10'd97;
assign feature_index_8[245] = 10'd655;
assign feature_index_8[246] = 10'd267;
assign feature_index_8[247] = 10'd348;
assign feature_index_8[248] = 10'd100;
assign feature_index_8[249] = 10'd441;
assign feature_index_8[250] = 10'd482;
assign feature_index_8[251] = 10'd314;
assign feature_index_8[252] = 10'd359;
assign feature_index_8[253] = 10'd343;
assign feature_index_8[254] = 10'd358;
assign feature_index_8[255] = 10'd371;
assign feature_index_8[256] = 10'd326;
assign feature_index_8[257] = 10'd400;
assign feature_index_8[258] = 10'd208;
assign feature_index_8[259] = 10'd436;
assign feature_index_8[260] = 10'd467;
assign feature_index_8[261] = 10'd491;
assign feature_index_8[262] = 10'd342;
assign feature_index_8[263] = 10'd581;
assign feature_index_8[264] = 10'd156;
assign feature_index_8[265] = 10'd490;
assign feature_index_8[266] = 10'd376;
assign feature_index_8[267] = 10'd405;
assign feature_index_8[268] = 10'd180;
assign feature_index_8[269] = 10'd520;
assign feature_index_8[270] = 10'd685;
assign feature_index_8[271] = 10'd712;
assign feature_index_8[272] = 10'd356;
assign feature_index_8[273] = 10'd569;
assign feature_index_8[274] = 10'd357;
assign feature_index_8[275] = 10'd401;
assign feature_index_8[276] = 10'd269;
assign feature_index_8[277] = 10'd377;
assign feature_index_8[278] = 10'd460;
assign feature_index_8[279] = 10'd430;
assign feature_index_8[280] = 10'd378;
assign feature_index_8[281] = 10'd387;
assign feature_index_8[282] = 10'd487;
assign feature_index_8[283] = 10'd686;
assign feature_index_8[284] = 10'd162;
assign feature_index_8[285] = 10'd426;
assign feature_index_8[286] = 10'd516;
assign feature_index_8[287] = 10'd566;
assign feature_index_8[288] = 10'd519;
assign feature_index_8[289] = 10'd154;
assign feature_index_8[290] = 10'd430;
assign feature_index_8[291] = 10'd154;
assign feature_index_8[292] = 10'd324;
assign feature_index_8[293] = 10'd319;
assign feature_index_8[294] = 10'd541;
assign feature_index_8[295] = 10'd428;
assign feature_index_8[296] = 10'd154;
assign feature_index_8[297] = 10'd207;
assign feature_index_8[298] = 10'd330;
assign feature_index_8[299] = 10'd416;
assign feature_index_8[300] = 10'd347;
assign feature_index_8[301] = 10'd121;
assign feature_index_8[302] = 10'd353;
assign feature_index_8[303] = 10'd684;
assign feature_index_8[304] = 10'd233;
assign feature_index_8[305] = 10'd575;
assign feature_index_8[306] = 10'd662;
assign feature_index_8[307] = 10'd0;
assign feature_index_8[308] = 10'd326;
assign feature_index_8[309] = 10'd405;
assign feature_index_8[310] = 10'd622;
assign feature_index_8[311] = 10'd375;
assign feature_index_8[312] = 10'd387;
assign feature_index_8[313] = 10'd298;
assign feature_index_8[314] = 10'd233;
assign feature_index_8[315] = 10'd493;
assign feature_index_8[316] = 10'd575;
assign feature_index_8[317] = 10'd488;
assign feature_index_8[318] = 10'd350;
assign feature_index_8[319] = 10'd266;
assign feature_index_8[320] = 10'd238;
assign feature_index_8[321] = 10'd180;
assign feature_index_8[322] = 10'd297;
assign feature_index_8[323] = 10'd397;
assign feature_index_8[324] = 10'd425;
assign feature_index_8[325] = 10'd356;
assign feature_index_8[326] = 10'd537;
assign feature_index_8[327] = 10'd651;
assign feature_index_8[328] = 10'd351;
assign feature_index_8[329] = 10'd545;
assign feature_index_8[330] = 10'd471;
assign feature_index_8[331] = 10'd489;
assign feature_index_8[332] = 10'd435;
assign feature_index_8[333] = 10'd630;
assign feature_index_8[334] = 10'd248;
assign feature_index_8[335] = 10'd181;
assign feature_index_8[336] = 10'd289;
assign feature_index_8[337] = 10'd316;
assign feature_index_8[338] = 10'd426;
assign feature_index_8[339] = 10'd227;
assign feature_index_8[340] = 10'd595;
assign feature_index_8[341] = 10'd341;
assign feature_index_8[342] = 10'd415;
assign feature_index_8[343] = 10'd294;
assign feature_index_8[344] = 10'd611;
assign feature_index_8[345] = 10'd0;
assign feature_index_8[346] = 10'd402;
assign feature_index_8[347] = 10'd344;
assign feature_index_8[348] = 10'd295;
assign feature_index_8[349] = 10'd183;
assign feature_index_8[350] = 10'd238;
assign feature_index_8[351] = 10'd182;
assign feature_index_8[352] = 10'd328;
assign feature_index_8[353] = 10'd271;
assign feature_index_8[354] = 10'd157;
assign feature_index_8[355] = 10'd544;
assign feature_index_8[356] = 10'd409;
assign feature_index_8[357] = 10'd237;
assign feature_index_8[358] = 10'd298;
assign feature_index_8[359] = 10'd381;
assign feature_index_8[360] = 10'd379;
assign feature_index_8[361] = 10'd264;
assign feature_index_8[362] = 10'd157;
assign feature_index_8[363] = 10'd161;
assign feature_index_8[364] = 10'd274;
assign feature_index_8[365] = 10'd569;
assign feature_index_8[366] = 10'd467;
assign feature_index_8[367] = 10'd331;
assign feature_index_8[368] = 10'd368;
assign feature_index_8[369] = 10'd189;
assign feature_index_8[370] = 10'd596;
assign feature_index_8[371] = 10'd162;
assign feature_index_8[372] = 10'd597;
assign feature_index_8[373] = 10'd0;
assign feature_index_8[374] = 10'd387;
assign feature_index_8[375] = 10'd655;
assign feature_index_8[376] = 10'd659;
assign feature_index_8[377] = 10'd486;
assign feature_index_8[378] = 10'd490;
assign feature_index_8[379] = 10'd244;
assign feature_index_8[380] = 10'd379;
assign feature_index_8[381] = 10'd432;
assign feature_index_8[382] = 10'd407;
assign feature_index_8[383] = 10'd271;
assign feature_index_8[384] = 10'd526;
assign feature_index_8[385] = 10'd352;
assign feature_index_8[386] = 10'd262;
assign feature_index_8[387] = 10'd683;
assign feature_index_8[388] = 10'd360;
assign feature_index_8[389] = 10'd658;
assign feature_index_8[390] = 10'd98;
assign feature_index_8[391] = 10'd626;
assign feature_index_8[392] = 10'd555;
assign feature_index_8[393] = 10'd0;
assign feature_index_8[394] = 10'd0;
assign feature_index_8[395] = 10'd0;
assign feature_index_8[396] = 10'd436;
assign feature_index_8[397] = 10'd0;
assign feature_index_8[398] = 10'd549;
assign feature_index_8[399] = 10'd539;
assign feature_index_8[400] = 10'd555;
assign feature_index_8[401] = 10'd206;
assign feature_index_8[402] = 10'd291;
assign feature_index_8[403] = 10'd551;
assign feature_index_8[404] = 10'd320;
assign feature_index_8[405] = 10'd381;
assign feature_index_8[406] = 10'd302;
assign feature_index_8[407] = 10'd516;
assign feature_index_8[408] = 10'd518;
assign feature_index_8[409] = 10'd187;
assign feature_index_8[410] = 10'd552;
assign feature_index_8[411] = 10'd161;
assign feature_index_8[412] = 10'd483;
assign feature_index_8[413] = 10'd189;
assign feature_index_8[414] = 10'd163;
assign feature_index_8[415] = 10'd302;
assign feature_index_8[416] = 10'd487;
assign feature_index_8[417] = 10'd328;
assign feature_index_8[418] = 10'd176;
assign feature_index_8[419] = 10'd414;
assign feature_index_8[420] = 10'd347;
assign feature_index_8[421] = 10'd347;
assign feature_index_8[422] = 10'd156;
assign feature_index_8[423] = 10'd486;
assign feature_index_8[424] = 10'd296;
assign feature_index_8[425] = 10'd712;
assign feature_index_8[426] = 10'd400;
assign feature_index_8[427] = 10'd626;
assign feature_index_8[428] = 10'd625;
assign feature_index_8[429] = 10'd297;
assign feature_index_8[430] = 10'd462;
assign feature_index_8[431] = 10'd354;
assign feature_index_8[432] = 10'd275;
assign feature_index_8[433] = 10'd542;
assign feature_index_8[434] = 10'd298;
assign feature_index_8[435] = 10'd345;
assign feature_index_8[436] = 10'd303;
assign feature_index_8[437] = 10'd711;
assign feature_index_8[438] = 10'd241;
assign feature_index_8[439] = 10'd583;
assign feature_index_8[440] = 10'd551;
assign feature_index_8[441] = 10'd327;
assign feature_index_8[442] = 10'd316;
assign feature_index_8[443] = 10'd219;
assign feature_index_8[444] = 10'd318;
assign feature_index_8[445] = 10'd272;
assign feature_index_8[446] = 10'd407;
assign feature_index_8[447] = 10'd427;
assign feature_index_8[448] = 10'd594;
assign feature_index_8[449] = 10'd0;
assign feature_index_8[450] = 10'd435;
assign feature_index_8[451] = 10'd178;
assign feature_index_8[452] = 10'd324;
assign feature_index_8[453] = 10'd383;
assign feature_index_8[454] = 10'd521;
assign feature_index_8[455] = 10'd297;
assign feature_index_8[456] = 10'd499;
assign feature_index_8[457] = 10'd0;
assign feature_index_8[458] = 10'd0;
assign feature_index_8[459] = 10'd161;
assign feature_index_8[460] = 10'd568;
assign feature_index_8[461] = 10'd527;
assign feature_index_8[462] = 10'd509;
assign feature_index_8[463] = 10'd714;
assign feature_index_8[464] = 10'd662;
assign feature_index_8[465] = 10'd595;
assign feature_index_8[466] = 10'd399;
assign feature_index_8[467] = 10'd383;
assign feature_index_8[468] = 10'd399;
assign feature_index_8[469] = 10'd460;
assign feature_index_8[470] = 10'd468;
assign feature_index_8[471] = 10'd515;
assign feature_index_8[472] = 10'd293;
assign feature_index_8[473] = 10'd0;
assign feature_index_8[474] = 10'd653;
assign feature_index_8[475] = 10'd299;
assign feature_index_8[476] = 10'd495;
assign feature_index_8[477] = 10'd461;
assign feature_index_8[478] = 10'd453;
assign feature_index_8[479] = 10'd380;
assign feature_index_8[480] = 10'd556;
assign feature_index_8[481] = 10'd581;
assign feature_index_8[482] = 10'd352;
assign feature_index_8[483] = 10'd499;
assign feature_index_8[484] = 10'd580;
assign feature_index_8[485] = 10'd470;
assign feature_index_8[486] = 10'd0;
assign feature_index_8[487] = 10'd246;
assign feature_index_8[488] = 10'd243;
assign feature_index_8[489] = 10'd691;
assign feature_index_8[490] = 10'd469;
assign feature_index_8[491] = 10'd576;
assign feature_index_8[492] = 10'd410;
assign feature_index_8[493] = 10'd482;
assign feature_index_8[494] = 10'd273;
assign feature_index_8[495] = 10'd359;
assign feature_index_8[496] = 10'd359;
assign feature_index_8[497] = 10'd149;
assign feature_index_8[498] = 10'd286;
assign feature_index_8[499] = 10'd344;
assign feature_index_8[500] = 10'd594;
assign feature_index_8[501] = 10'd431;
assign feature_index_8[502] = 10'd154;
assign feature_index_8[503] = 10'd316;
assign feature_index_8[504] = 10'd370;
assign feature_index_8[505] = 10'd523;
assign feature_index_8[506] = 10'd260;
assign feature_index_8[507] = 10'd660;
assign feature_index_8[508] = 10'd601;
assign feature_index_8[509] = 10'd185;
assign feature_index_8[510] = 10'd468;
assign feature_index_8[511] = 10'd128;
assign feature_index_8[512] = 10'd183;
assign feature_index_8[513] = 10'd219;
assign feature_index_8[514] = 10'd406;
assign feature_index_8[515] = 10'd297;
assign feature_index_8[516] = 10'd325;
assign feature_index_8[517] = 10'd655;
assign feature_index_8[518] = 10'd405;
assign feature_index_8[519] = 10'd151;
assign feature_index_8[520] = 10'd377;
assign feature_index_8[521] = 10'd469;
assign feature_index_8[522] = 10'd405;
assign feature_index_8[523] = 10'd149;
assign feature_index_8[524] = 10'd358;
assign feature_index_8[525] = 10'd0;
assign feature_index_8[526] = 10'd179;
assign feature_index_8[527] = 10'd539;
assign feature_index_8[528] = 10'd320;
assign feature_index_8[529] = 10'd487;
assign feature_index_8[530] = 10'd375;
assign feature_index_8[531] = 10'd276;
assign feature_index_8[532] = 10'd712;
assign feature_index_8[533] = 10'd526;
assign feature_index_8[534] = 10'd324;
assign feature_index_8[535] = 10'd567;
assign feature_index_8[536] = 10'd627;
assign feature_index_8[537] = 10'd208;
assign feature_index_8[538] = 10'd125;
assign feature_index_8[539] = 10'd330;
assign feature_index_8[540] = 10'd323;
assign feature_index_8[541] = 10'd341;
assign feature_index_8[542] = 10'd343;
assign feature_index_8[543] = 10'd536;
assign feature_index_8[544] = 10'd0;
assign feature_index_8[545] = 10'd710;
assign feature_index_8[546] = 10'd301;
assign feature_index_8[547] = 10'd486;
assign feature_index_8[548] = 10'd352;
assign feature_index_8[549] = 10'd602;
assign feature_index_8[550] = 10'd159;
assign feature_index_8[551] = 10'd563;
assign feature_index_8[552] = 10'd378;
assign feature_index_8[553] = 10'd271;
assign feature_index_8[554] = 10'd0;
assign feature_index_8[555] = 10'd488;
assign feature_index_8[556] = 10'd185;
assign feature_index_8[557] = 10'd211;
assign feature_index_8[558] = 10'd655;
assign feature_index_8[559] = 10'd410;
assign feature_index_8[560] = 10'd487;
assign feature_index_8[561] = 10'd371;
assign feature_index_8[562] = 10'd373;
assign feature_index_8[563] = 10'd683;
assign feature_index_8[564] = 10'd0;
assign feature_index_8[565] = 10'd153;
assign feature_index_8[566] = 10'd156;
assign feature_index_8[567] = 10'd405;
assign feature_index_8[568] = 10'd689;
assign feature_index_8[569] = 10'd0;
assign feature_index_8[570] = 10'd0;
assign feature_index_8[571] = 10'd599;
assign feature_index_8[572] = 10'd465;
assign feature_index_8[573] = 10'd521;
assign feature_index_8[574] = 10'd434;
assign feature_index_8[575] = 10'd348;
assign feature_index_8[576] = 10'd490;
assign feature_index_8[577] = 10'd317;
assign feature_index_8[578] = 10'd405;
assign feature_index_8[579] = 10'd536;
assign feature_index_8[580] = 10'd318;
assign feature_index_8[581] = 10'd598;
assign feature_index_8[582] = 10'd455;
assign feature_index_8[583] = 10'd552;
assign feature_index_8[584] = 10'd424;
assign feature_index_8[585] = 10'd319;
assign feature_index_8[586] = 10'd263;
assign feature_index_8[587] = 10'd711;
assign feature_index_8[588] = 10'd295;
assign feature_index_8[589] = 10'd379;
assign feature_index_8[590] = 10'd97;
assign feature_index_8[591] = 10'd377;
assign feature_index_8[592] = 10'd377;
assign feature_index_8[593] = 10'd713;
assign feature_index_8[594] = 10'd545;
assign feature_index_8[595] = 10'd208;
assign feature_index_8[596] = 10'd628;
assign feature_index_8[597] = 10'd152;
assign feature_index_8[598] = 10'd510;
assign feature_index_8[599] = 10'd605;
assign feature_index_8[600] = 10'd0;
assign feature_index_8[601] = 10'd523;
assign feature_index_8[602] = 10'd0;
assign feature_index_8[603] = 10'd379;
assign feature_index_8[604] = 10'd0;
assign feature_index_8[605] = 10'd0;
assign feature_index_8[606] = 10'd464;
assign feature_index_8[607] = 10'd547;
assign feature_index_8[608] = 10'd319;
assign feature_index_8[609] = 10'd656;
assign feature_index_8[610] = 10'd239;
assign feature_index_8[611] = 10'd541;
assign feature_index_8[612] = 10'd264;
assign feature_index_8[613] = 10'd270;
assign feature_index_8[614] = 10'd120;
assign feature_index_8[615] = 10'd0;
assign feature_index_8[616] = 10'd0;
assign feature_index_8[617] = 10'd0;
assign feature_index_8[618] = 10'd0;
assign feature_index_8[619] = 10'd689;
assign feature_index_8[620] = 10'd178;
assign feature_index_8[621] = 10'd570;
assign feature_index_8[622] = 10'd406;
assign feature_index_8[623] = 10'd544;
assign feature_index_8[624] = 10'd578;
assign feature_index_8[625] = 10'd377;
assign feature_index_8[626] = 10'd215;
assign feature_index_8[627] = 10'd101;
assign feature_index_8[628] = 10'd404;
assign feature_index_8[629] = 10'd430;
assign feature_index_8[630] = 10'd321;
assign feature_index_8[631] = 10'd516;
assign feature_index_8[632] = 10'd595;
assign feature_index_8[633] = 10'd329;
assign feature_index_8[634] = 10'd488;
assign feature_index_8[635] = 10'd347;
assign feature_index_8[636] = 10'd666;
assign feature_index_8[637] = 10'd466;
assign feature_index_8[638] = 10'd0;
assign feature_index_8[639] = 10'd514;
assign feature_index_8[640] = 10'd430;
assign feature_index_8[641] = 10'd182;
assign feature_index_8[642] = 10'd432;
assign feature_index_8[643] = 10'd178;
assign feature_index_8[644] = 10'd437;
assign feature_index_8[645] = 10'd377;
assign feature_index_8[646] = 10'd376;
assign feature_index_8[647] = 10'd130;
assign feature_index_8[648] = 10'd266;
assign feature_index_8[649] = 10'd496;
assign feature_index_8[650] = 10'd271;
assign feature_index_8[651] = 10'd0;
assign feature_index_8[652] = 10'd408;
assign feature_index_8[653] = 10'd0;
assign feature_index_8[654] = 10'd276;
assign feature_index_8[655] = 10'd292;
assign feature_index_8[656] = 10'd630;
assign feature_index_8[657] = 10'd403;
assign feature_index_8[658] = 10'd204;
assign feature_index_8[659] = 10'd544;
assign feature_index_8[660] = 10'd659;
assign feature_index_8[661] = 10'd411;
assign feature_index_8[662] = 10'd291;
assign feature_index_8[663] = 10'd358;
assign feature_index_8[664] = 10'd356;
assign feature_index_8[665] = 10'd415;
assign feature_index_8[666] = 10'd248;
assign feature_index_8[667] = 10'd579;
assign feature_index_8[668] = 10'd516;
assign feature_index_8[669] = 10'd263;
assign feature_index_8[670] = 10'd128;
assign feature_index_8[671] = 10'd565;
assign feature_index_8[672] = 10'd536;
assign feature_index_8[673] = 10'd294;
assign feature_index_8[674] = 10'd487;
assign feature_index_8[675] = 10'd323;
assign feature_index_8[676] = 10'd452;
assign feature_index_8[677] = 10'd302;
assign feature_index_8[678] = 10'd409;
assign feature_index_8[679] = 10'd269;
assign feature_index_8[680] = 10'd0;
assign feature_index_8[681] = 10'd655;
assign feature_index_8[682] = 10'd398;
assign feature_index_8[683] = 10'd376;
assign feature_index_8[684] = 10'd406;
assign feature_index_8[685] = 10'd359;
assign feature_index_8[686] = 10'd427;
assign feature_index_8[687] = 10'd273;
assign feature_index_8[688] = 10'd175;
assign feature_index_8[689] = 10'd0;
assign feature_index_8[690] = 10'd184;
assign feature_index_8[691] = 10'd0;
assign feature_index_8[692] = 10'd0;
assign feature_index_8[693] = 10'd0;
assign feature_index_8[694] = 10'd0;
assign feature_index_8[695] = 10'd126;
assign feature_index_8[696] = 10'd233;
assign feature_index_8[697] = 10'd355;
assign feature_index_8[698] = 10'd289;
assign feature_index_8[699] = 10'd400;
assign feature_index_8[700] = 10'd228;
assign feature_index_8[701] = 10'd0;
assign feature_index_8[702] = 10'd386;
assign feature_index_8[703] = 10'd96;
assign feature_index_8[704] = 10'd467;
assign feature_index_8[705] = 10'd160;
assign feature_index_8[706] = 10'd220;
assign feature_index_8[707] = 10'd231;
assign feature_index_8[708] = 10'd261;
assign feature_index_8[709] = 10'd274;
assign feature_index_8[710] = 10'd632;
assign feature_index_8[711] = 10'd497;
assign feature_index_8[712] = 10'd711;
assign feature_index_8[713] = 10'd608;
assign feature_index_8[714] = 10'd579;
assign feature_index_8[715] = 10'd608;
assign feature_index_8[716] = 10'd552;
assign feature_index_8[717] = 10'd318;
assign feature_index_8[718] = 10'd412;
assign feature_index_8[719] = 10'd454;
assign feature_index_8[720] = 10'd130;
assign feature_index_8[721] = 10'd382;
assign feature_index_8[722] = 10'd659;
assign feature_index_8[723] = 10'd263;
assign feature_index_8[724] = 10'd234;
assign feature_index_8[725] = 10'd464;
assign feature_index_8[726] = 10'd294;
assign feature_index_8[727] = 10'd249;
assign feature_index_8[728] = 10'd192;
assign feature_index_8[729] = 10'd295;
assign feature_index_8[730] = 10'd538;
assign feature_index_8[731] = 10'd160;
assign feature_index_8[732] = 10'd185;
assign feature_index_8[733] = 10'd660;
assign feature_index_8[734] = 10'd624;
assign feature_index_8[735] = 10'd264;
assign feature_index_8[736] = 10'd0;
assign feature_index_8[737] = 10'd623;
assign feature_index_8[738] = 10'd0;
assign feature_index_8[739] = 10'd0;
assign feature_index_8[740] = 10'd572;
assign feature_index_8[741] = 10'd180;
assign feature_index_8[742] = 10'd0;
assign feature_index_8[743] = 10'd387;
assign feature_index_8[744] = 10'd315;
assign feature_index_8[745] = 10'd404;
assign feature_index_8[746] = 10'd236;
assign feature_index_8[747] = 10'd0;
assign feature_index_8[748] = 10'd0;
assign feature_index_8[749] = 10'd149;
assign feature_index_8[750] = 10'd238;
assign feature_index_8[751] = 10'd183;
assign feature_index_8[752] = 10'd380;
assign feature_index_8[753] = 10'd244;
assign feature_index_8[754] = 10'd243;
assign feature_index_8[755] = 10'd0;
assign feature_index_8[756] = 10'd267;
assign feature_index_8[757] = 10'd350;
assign feature_index_8[758] = 10'd186;
assign feature_index_8[759] = 10'd628;
assign feature_index_8[760] = 10'd353;
assign feature_index_8[761] = 10'd298;
assign feature_index_8[762] = 10'd657;
assign feature_index_8[763] = 10'd270;
assign feature_index_8[764] = 10'd542;
assign feature_index_8[765] = 10'd275;
assign feature_index_8[766] = 10'd182;
assign feature_index_8[767] = 10'd383;
assign feature_index_8[768] = 10'd402;
assign feature_index_8[769] = 10'd471;
assign feature_index_8[770] = 10'd608;
assign feature_index_8[771] = 10'd432;
assign feature_index_8[772] = 10'd211;
assign feature_index_8[773] = 10'd259;
assign feature_index_8[774] = 10'd237;
assign feature_index_8[775] = 10'd600;
assign feature_index_8[776] = 10'd601;
assign feature_index_8[777] = 10'd184;
assign feature_index_8[778] = 10'd0;
assign feature_index_8[779] = 10'd294;
assign feature_index_8[780] = 10'd0;
assign feature_index_8[781] = 10'd492;
assign feature_index_8[782] = 10'd0;
assign feature_index_8[783] = 10'd0;
assign feature_index_8[784] = 10'd544;
assign feature_index_8[785] = 10'd0;
assign feature_index_8[786] = 10'd0;
assign feature_index_8[787] = 10'd0;
assign feature_index_8[788] = 10'd0;
assign feature_index_8[789] = 10'd0;
assign feature_index_8[790] = 10'd0;
assign feature_index_8[791] = 10'd0;
assign feature_index_8[792] = 10'd0;
assign feature_index_8[793] = 10'd354;
assign feature_index_8[794] = 10'd0;
assign feature_index_8[795] = 10'd0;
assign feature_index_8[796] = 10'd0;
assign feature_index_8[797] = 10'd0;
assign feature_index_8[798] = 10'd0;
assign feature_index_8[799] = 10'd209;
assign feature_index_8[800] = 10'd454;
assign feature_index_8[801] = 10'd370;
assign feature_index_8[802] = 10'd453;
assign feature_index_8[803] = 10'd500;
assign feature_index_8[804] = 10'd318;
assign feature_index_8[805] = 10'd127;
assign feature_index_8[806] = 10'd240;
assign feature_index_8[807] = 10'd217;
assign feature_index_8[808] = 10'd386;
assign feature_index_8[809] = 10'd100;
assign feature_index_8[810] = 10'd571;
assign feature_index_8[811] = 10'd0;
assign feature_index_8[812] = 10'd621;
assign feature_index_8[813] = 10'd260;
assign feature_index_8[814] = 10'd210;
assign feature_index_8[815] = 10'd520;
assign feature_index_8[816] = 10'd0;
assign feature_index_8[817] = 10'd0;
assign feature_index_8[818] = 10'd173;
assign feature_index_8[819] = 10'd236;
assign feature_index_8[820] = 10'd405;
assign feature_index_8[821] = 10'd210;
assign feature_index_8[822] = 10'd0;
assign feature_index_8[823] = 10'd0;
assign feature_index_8[824] = 10'd0;
assign feature_index_8[825] = 10'd569;
assign feature_index_8[826] = 10'd538;
assign feature_index_8[827] = 10'd512;
assign feature_index_8[828] = 10'd156;
assign feature_index_8[829] = 10'd299;
assign feature_index_8[830] = 10'd0;
assign feature_index_8[831] = 10'd436;
assign feature_index_8[832] = 10'd567;
assign feature_index_8[833] = 10'd0;
assign feature_index_8[834] = 10'd185;
assign feature_index_8[835] = 10'd326;
assign feature_index_8[836] = 10'd400;
assign feature_index_8[837] = 10'd329;
assign feature_index_8[838] = 10'd288;
assign feature_index_8[839] = 10'd407;
assign feature_index_8[840] = 10'd0;
assign feature_index_8[841] = 10'd631;
assign feature_index_8[842] = 10'd655;
assign feature_index_8[843] = 10'd263;
assign feature_index_8[844] = 10'd0;
assign feature_index_8[845] = 10'd357;
assign feature_index_8[846] = 10'd495;
assign feature_index_8[847] = 10'd538;
assign feature_index_8[848] = 10'd348;
assign feature_index_8[849] = 10'd397;
assign feature_index_8[850] = 10'd466;
assign feature_index_8[851] = 10'd463;
assign feature_index_8[852] = 10'd242;
assign feature_index_8[853] = 10'd0;
assign feature_index_8[854] = 10'd410;
assign feature_index_8[855] = 10'd711;
assign feature_index_8[856] = 10'd548;
assign feature_index_8[857] = 10'd273;
assign feature_index_8[858] = 10'd377;
assign feature_index_8[859] = 10'd578;
assign feature_index_8[860] = 10'd212;
assign feature_index_8[861] = 10'd380;
assign feature_index_8[862] = 10'd192;
assign feature_index_8[863] = 10'd598;
assign feature_index_8[864] = 10'd521;
assign feature_index_8[865] = 10'd131;
assign feature_index_8[866] = 10'd401;
assign feature_index_8[867] = 10'd512;
assign feature_index_8[868] = 10'd512;
assign feature_index_8[869] = 10'd383;
assign feature_index_8[870] = 10'd539;
assign feature_index_8[871] = 10'd370;
assign feature_index_8[872] = 10'd257;
assign feature_index_8[873] = 10'd372;
assign feature_index_8[874] = 10'd497;
assign feature_index_8[875] = 10'd577;
assign feature_index_8[876] = 10'd247;
assign feature_index_8[877] = 10'd596;
assign feature_index_8[878] = 10'd485;
assign feature_index_8[879] = 10'd636;
assign feature_index_8[880] = 10'd0;
assign feature_index_8[881] = 10'd542;
assign feature_index_8[882] = 10'd461;
assign feature_index_8[883] = 10'd269;
assign feature_index_8[884] = 10'd657;
assign feature_index_8[885] = 10'd156;
assign feature_index_8[886] = 10'd402;
assign feature_index_8[887] = 10'd268;
assign feature_index_8[888] = 10'd105;
assign feature_index_8[889] = 10'd296;
assign feature_index_8[890] = 10'd400;
assign feature_index_8[891] = 10'd373;
assign feature_index_8[892] = 10'd123;
assign feature_index_8[893] = 10'd520;
assign feature_index_8[894] = 10'd297;
assign feature_index_8[895] = 10'd318;
assign feature_index_8[896] = 10'd566;
assign feature_index_8[897] = 10'd258;
assign feature_index_8[898] = 10'd160;
assign feature_index_8[899] = 10'd0;
assign feature_index_8[900] = 10'd0;
assign feature_index_8[901] = 10'd0;
assign feature_index_8[902] = 10'd0;
assign feature_index_8[903] = 10'd0;
assign feature_index_8[904] = 10'd438;
assign feature_index_8[905] = 10'd192;
assign feature_index_8[906] = 10'd0;
assign feature_index_8[907] = 10'd131;
assign feature_index_8[908] = 10'd638;
assign feature_index_8[909] = 10'd127;
assign feature_index_8[910] = 10'd564;
assign feature_index_8[911] = 10'd593;
assign feature_index_8[912] = 10'd346;
assign feature_index_8[913] = 10'd512;
assign feature_index_8[914] = 10'd0;
assign feature_index_8[915] = 10'd0;
assign feature_index_8[916] = 10'd0;
assign feature_index_8[917] = 10'd0;
assign feature_index_8[918] = 10'd0;
assign feature_index_8[919] = 10'd0;
assign feature_index_8[920] = 10'd607;
assign feature_index_8[921] = 10'd0;
assign feature_index_8[922] = 10'd248;
assign feature_index_8[923] = 10'd0;
assign feature_index_8[924] = 10'd127;
assign feature_index_8[925] = 10'd0;
assign feature_index_8[926] = 10'd0;
assign feature_index_8[927] = 10'd288;
assign feature_index_8[928] = 10'd459;
assign feature_index_8[929] = 10'd153;
assign feature_index_8[930] = 10'd0;
assign feature_index_8[931] = 10'd245;
assign feature_index_8[932] = 10'd273;
assign feature_index_8[933] = 10'd624;
assign feature_index_8[934] = 10'd0;
assign feature_index_8[935] = 10'd463;
assign feature_index_8[936] = 10'd522;
assign feature_index_8[937] = 10'd598;
assign feature_index_8[938] = 10'd571;
assign feature_index_8[939] = 10'd0;
assign feature_index_8[940] = 10'd274;
assign feature_index_8[941] = 10'd0;
assign feature_index_8[942] = 10'd0;
assign feature_index_8[943] = 10'd497;
assign feature_index_8[944] = 10'd136;
assign feature_index_8[945] = 10'd378;
assign feature_index_8[946] = 10'd303;
assign feature_index_8[947] = 10'd0;
assign feature_index_8[948] = 10'd0;
assign feature_index_8[949] = 10'd516;
assign feature_index_8[950] = 10'd0;
assign feature_index_8[951] = 10'd193;
assign feature_index_8[952] = 10'd408;
assign feature_index_8[953] = 10'd206;
assign feature_index_8[954] = 10'd0;
assign feature_index_8[955] = 10'd237;
assign feature_index_8[956] = 10'd599;
assign feature_index_8[957] = 10'd399;
assign feature_index_8[958] = 10'd0;
assign feature_index_8[959] = 10'd126;
assign feature_index_8[960] = 10'd606;
assign feature_index_8[961] = 10'd181;
assign feature_index_8[962] = 10'd0;
assign feature_index_8[963] = 10'd499;
assign feature_index_8[964] = 10'd574;
assign feature_index_8[965] = 10'd289;
assign feature_index_8[966] = 10'd517;
assign feature_index_8[967] = 10'd383;
assign feature_index_8[968] = 10'd120;
assign feature_index_8[969] = 10'd541;
assign feature_index_8[970] = 10'd0;
assign feature_index_8[971] = 10'd217;
assign feature_index_8[972] = 10'd666;
assign feature_index_8[973] = 10'd0;
assign feature_index_8[974] = 10'd0;
assign feature_index_8[975] = 10'd155;
assign feature_index_8[976] = 10'd551;
assign feature_index_8[977] = 10'd341;
assign feature_index_8[978] = 10'd93;
assign feature_index_8[979] = 10'd72;
assign feature_index_8[980] = 10'd599;
assign feature_index_8[981] = 10'd537;
assign feature_index_8[982] = 10'd0;
assign feature_index_8[983] = 10'd245;
assign feature_index_8[984] = 10'd187;
assign feature_index_8[985] = 10'd0;
assign feature_index_8[986] = 10'd622;
assign feature_index_8[987] = 10'd537;
assign feature_index_8[988] = 10'd0;
assign feature_index_8[989] = 10'd682;
assign feature_index_8[990] = 10'd159;
assign feature_index_8[991] = 10'd471;
assign feature_index_8[992] = 10'd323;
assign feature_index_8[993] = 10'd123;
assign feature_index_8[994] = 10'd0;
assign feature_index_8[995] = 10'd567;
assign feature_index_8[996] = 10'd351;
assign feature_index_8[997] = 10'd0;
assign feature_index_8[998] = 10'd0;
assign feature_index_8[999] = 10'd719;
assign feature_index_8[1000] = 10'd219;
assign feature_index_8[1001] = 10'd344;
assign feature_index_8[1002] = 10'd0;
assign feature_index_8[1003] = 10'd630;
assign feature_index_8[1004] = 10'd681;
assign feature_index_8[1005] = 10'd634;
assign feature_index_8[1006] = 10'd579;
assign feature_index_8[1007] = 10'd681;
assign feature_index_8[1008] = 10'd399;
assign feature_index_8[1009] = 10'd470;
assign feature_index_8[1010] = 10'd94;
assign feature_index_8[1011] = 10'd626;
assign feature_index_8[1012] = 10'd526;
assign feature_index_8[1013] = 10'd0;
assign feature_index_8[1014] = 10'd0;
assign feature_index_8[1015] = 10'd319;
assign feature_index_8[1016] = 10'd580;
assign feature_index_8[1017] = 10'd403;
assign feature_index_8[1018] = 10'd545;
assign feature_index_8[1019] = 10'd295;
assign feature_index_8[1020] = 10'd462;
assign feature_index_8[1021] = 10'd515;
assign feature_index_8[1022] = 10'd267;
assign feature_index_9[0] = 10'd462;
assign feature_index_9[1] = 10'd301;
assign feature_index_9[2] = 10'd569;
assign feature_index_9[3] = 10'd628;
assign feature_index_9[4] = 10'd455;
assign feature_index_9[5] = 10'd428;
assign feature_index_9[6] = 10'd127;
assign feature_index_9[7] = 10'd742;
assign feature_index_9[8] = 10'd289;
assign feature_index_9[9] = 10'd156;
assign feature_index_9[10] = 10'd599;
assign feature_index_9[11] = 10'd318;
assign feature_index_9[12] = 10'd209;
assign feature_index_9[13] = 10'd182;
assign feature_index_9[14] = 10'd269;
assign feature_index_9[15] = 10'd326;
assign feature_index_9[16] = 10'd377;
assign feature_index_9[17] = 10'd295;
assign feature_index_9[18] = 10'd711;
assign feature_index_9[19] = 10'd411;
assign feature_index_9[20] = 10'd380;
assign feature_index_9[21] = 10'd180;
assign feature_index_9[22] = 10'd185;
assign feature_index_9[23] = 10'd244;
assign feature_index_9[24] = 10'd184;
assign feature_index_9[25] = 10'd709;
assign feature_index_9[26] = 10'd319;
assign feature_index_9[27] = 10'd247;
assign feature_index_9[28] = 10'd319;
assign feature_index_9[29] = 10'd513;
assign feature_index_9[30] = 10'd124;
assign feature_index_9[31] = 10'd98;
assign feature_index_9[32] = 10'd294;
assign feature_index_9[33] = 10'd233;
assign feature_index_9[34] = 10'd340;
assign feature_index_9[35] = 10'd351;
assign feature_index_9[36] = 10'd179;
assign feature_index_9[37] = 10'd360;
assign feature_index_9[38] = 10'd186;
assign feature_index_9[39] = 10'd524;
assign feature_index_9[40] = 10'd434;
assign feature_index_9[41] = 10'd622;
assign feature_index_9[42] = 10'd485;
assign feature_index_9[43] = 10'd567;
assign feature_index_9[44] = 10'd655;
assign feature_index_9[45] = 10'd409;
assign feature_index_9[46] = 10'd409;
assign feature_index_9[47] = 10'd458;
assign feature_index_9[48] = 10'd378;
assign feature_index_9[49] = 10'd267;
assign feature_index_9[50] = 10'd409;
assign feature_index_9[51] = 10'd98;
assign feature_index_9[52] = 10'd213;
assign feature_index_9[53] = 10'd378;
assign feature_index_9[54] = 10'd240;
assign feature_index_9[55] = 10'd548;
assign feature_index_9[56] = 10'd489;
assign feature_index_9[57] = 10'd657;
assign feature_index_9[58] = 10'd327;
assign feature_index_9[59] = 10'd595;
assign feature_index_9[60] = 10'd300;
assign feature_index_9[61] = 10'd350;
assign feature_index_9[62] = 10'd515;
assign feature_index_9[63] = 10'd101;
assign feature_index_9[64] = 10'd157;
assign feature_index_9[65] = 10'd125;
assign feature_index_9[66] = 10'd457;
assign feature_index_9[67] = 10'd487;
assign feature_index_9[68] = 10'd460;
assign feature_index_9[69] = 10'd413;
assign feature_index_9[70] = 10'd431;
assign feature_index_9[71] = 10'd518;
assign feature_index_9[72] = 10'd163;
assign feature_index_9[73] = 10'd456;
assign feature_index_9[74] = 10'd488;
assign feature_index_9[75] = 10'd349;
assign feature_index_9[76] = 10'd122;
assign feature_index_9[77] = 10'd318;
assign feature_index_9[78] = 10'd299;
assign feature_index_9[79] = 10'd353;
assign feature_index_9[80] = 10'd240;
assign feature_index_9[81] = 10'd593;
assign feature_index_9[82] = 10'd467;
assign feature_index_9[83] = 10'd276;
assign feature_index_9[84] = 10'd464;
assign feature_index_9[85] = 10'd595;
assign feature_index_9[86] = 10'd384;
assign feature_index_9[87] = 10'd213;
assign feature_index_9[88] = 10'd665;
assign feature_index_9[89] = 10'd498;
assign feature_index_9[90] = 10'd491;
assign feature_index_9[91] = 10'd459;
assign feature_index_9[92] = 10'd241;
assign feature_index_9[93] = 10'd563;
assign feature_index_9[94] = 10'd412;
assign feature_index_9[95] = 10'd203;
assign feature_index_9[96] = 10'd543;
assign feature_index_9[97] = 10'd458;
assign feature_index_9[98] = 10'd293;
assign feature_index_9[99] = 10'd153;
assign feature_index_9[100] = 10'd626;
assign feature_index_9[101] = 10'd517;
assign feature_index_9[102] = 10'd661;
assign feature_index_9[103] = 10'd67;
assign feature_index_9[104] = 10'd213;
assign feature_index_9[105] = 10'd289;
assign feature_index_9[106] = 10'd207;
assign feature_index_9[107] = 10'd409;
assign feature_index_9[108] = 10'd653;
assign feature_index_9[109] = 10'd552;
assign feature_index_9[110] = 10'd442;
assign feature_index_9[111] = 10'd400;
assign feature_index_9[112] = 10'd429;
assign feature_index_9[113] = 10'd329;
assign feature_index_9[114] = 10'd653;
assign feature_index_9[115] = 10'd652;
assign feature_index_9[116] = 10'd151;
assign feature_index_9[117] = 10'd410;
assign feature_index_9[118] = 10'd654;
assign feature_index_9[119] = 10'd383;
assign feature_index_9[120] = 10'd323;
assign feature_index_9[121] = 10'd656;
assign feature_index_9[122] = 10'd496;
assign feature_index_9[123] = 10'd293;
assign feature_index_9[124] = 10'd525;
assign feature_index_9[125] = 10'd378;
assign feature_index_9[126] = 10'd603;
assign feature_index_9[127] = 10'd218;
assign feature_index_9[128] = 10'd183;
assign feature_index_9[129] = 10'd246;
assign feature_index_9[130] = 10'd289;
assign feature_index_9[131] = 10'd239;
assign feature_index_9[132] = 10'd567;
assign feature_index_9[133] = 10'd186;
assign feature_index_9[134] = 10'd543;
assign feature_index_9[135] = 10'd406;
assign feature_index_9[136] = 10'd381;
assign feature_index_9[137] = 10'd402;
assign feature_index_9[138] = 10'd317;
assign feature_index_9[139] = 10'd404;
assign feature_index_9[140] = 10'd374;
assign feature_index_9[141] = 10'd0;
assign feature_index_9[142] = 10'd0;
assign feature_index_9[143] = 10'd405;
assign feature_index_9[144] = 10'd153;
assign feature_index_9[145] = 10'd299;
assign feature_index_9[146] = 10'd272;
assign feature_index_9[147] = 10'd246;
assign feature_index_9[148] = 10'd429;
assign feature_index_9[149] = 10'd378;
assign feature_index_9[150] = 10'd528;
assign feature_index_9[151] = 10'd408;
assign feature_index_9[152] = 10'd487;
assign feature_index_9[153] = 10'd149;
assign feature_index_9[154] = 10'd347;
assign feature_index_9[155] = 10'd376;
assign feature_index_9[156] = 10'd430;
assign feature_index_9[157] = 10'd354;
assign feature_index_9[158] = 10'd518;
assign feature_index_9[159] = 10'd442;
assign feature_index_9[160] = 10'd321;
assign feature_index_9[161] = 10'd713;
assign feature_index_9[162] = 10'd436;
assign feature_index_9[163] = 10'd405;
assign feature_index_9[164] = 10'd349;
assign feature_index_9[165] = 10'd594;
assign feature_index_9[166] = 10'd653;
assign feature_index_9[167] = 10'd538;
assign feature_index_9[168] = 10'd495;
assign feature_index_9[169] = 10'd353;
assign feature_index_9[170] = 10'd375;
assign feature_index_9[171] = 10'd290;
assign feature_index_9[172] = 10'd289;
assign feature_index_9[173] = 10'd317;
assign feature_index_9[174] = 10'd322;
assign feature_index_9[175] = 10'd543;
assign feature_index_9[176] = 10'd434;
assign feature_index_9[177] = 10'd239;
assign feature_index_9[178] = 10'd270;
assign feature_index_9[179] = 10'd428;
assign feature_index_9[180] = 10'd415;
assign feature_index_9[181] = 10'd381;
assign feature_index_9[182] = 10'd267;
assign feature_index_9[183] = 10'd325;
assign feature_index_9[184] = 10'd131;
assign feature_index_9[185] = 10'd495;
assign feature_index_9[186] = 10'd329;
assign feature_index_9[187] = 10'd408;
assign feature_index_9[188] = 10'd154;
assign feature_index_9[189] = 10'd598;
assign feature_index_9[190] = 10'd265;
assign feature_index_9[191] = 10'd262;
assign feature_index_9[192] = 10'd519;
assign feature_index_9[193] = 10'd546;
assign feature_index_9[194] = 10'd324;
assign feature_index_9[195] = 10'd354;
assign feature_index_9[196] = 10'd157;
assign feature_index_9[197] = 10'd543;
assign feature_index_9[198] = 10'd221;
assign feature_index_9[199] = 10'd469;
assign feature_index_9[200] = 10'd98;
assign feature_index_9[201] = 10'd230;
assign feature_index_9[202] = 10'd383;
assign feature_index_9[203] = 10'd352;
assign feature_index_9[204] = 10'd543;
assign feature_index_9[205] = 10'd155;
assign feature_index_9[206] = 10'd542;
assign feature_index_9[207] = 10'd266;
assign feature_index_9[208] = 10'd0;
assign feature_index_9[209] = 10'd481;
assign feature_index_9[210] = 10'd0;
assign feature_index_9[211] = 10'd461;
assign feature_index_9[212] = 10'd240;
assign feature_index_9[213] = 10'd459;
assign feature_index_9[214] = 10'd629;
assign feature_index_9[215] = 10'd481;
assign feature_index_9[216] = 10'd151;
assign feature_index_9[217] = 10'd318;
assign feature_index_9[218] = 10'd605;
assign feature_index_9[219] = 10'd186;
assign feature_index_9[220] = 10'd691;
assign feature_index_9[221] = 10'd193;
assign feature_index_9[222] = 10'd201;
assign feature_index_9[223] = 10'd378;
assign feature_index_9[224] = 10'd95;
assign feature_index_9[225] = 10'd656;
assign feature_index_9[226] = 10'd572;
assign feature_index_9[227] = 10'd326;
assign feature_index_9[228] = 10'd162;
assign feature_index_9[229] = 10'd410;
assign feature_index_9[230] = 10'd411;
assign feature_index_9[231] = 10'd370;
assign feature_index_9[232] = 10'd550;
assign feature_index_9[233] = 10'd550;
assign feature_index_9[234] = 10'd429;
assign feature_index_9[235] = 10'd245;
assign feature_index_9[236] = 10'd658;
assign feature_index_9[237] = 10'd74;
assign feature_index_9[238] = 10'd684;
assign feature_index_9[239] = 10'd270;
assign feature_index_9[240] = 10'd568;
assign feature_index_9[241] = 10'd158;
assign feature_index_9[242] = 10'd299;
assign feature_index_9[243] = 10'd216;
assign feature_index_9[244] = 10'd354;
assign feature_index_9[245] = 10'd324;
assign feature_index_9[246] = 10'd187;
assign feature_index_9[247] = 10'd344;
assign feature_index_9[248] = 10'd326;
assign feature_index_9[249] = 10'd576;
assign feature_index_9[250] = 10'd316;
assign feature_index_9[251] = 10'd381;
assign feature_index_9[252] = 10'd458;
assign feature_index_9[253] = 10'd627;
assign feature_index_9[254] = 10'd347;
assign feature_index_9[255] = 10'd545;
assign feature_index_9[256] = 10'd381;
assign feature_index_9[257] = 10'd600;
assign feature_index_9[258] = 10'd296;
assign feature_index_9[259] = 10'd324;
assign feature_index_9[260] = 10'd578;
assign feature_index_9[261] = 10'd436;
assign feature_index_9[262] = 10'd596;
assign feature_index_9[263] = 10'd682;
assign feature_index_9[264] = 10'd230;
assign feature_index_9[265] = 10'd242;
assign feature_index_9[266] = 10'd387;
assign feature_index_9[267] = 10'd401;
assign feature_index_9[268] = 10'd268;
assign feature_index_9[269] = 10'd434;
assign feature_index_9[270] = 10'd242;
assign feature_index_9[271] = 10'd316;
assign feature_index_9[272] = 10'd0;
assign feature_index_9[273] = 10'd0;
assign feature_index_9[274] = 10'd0;
assign feature_index_9[275] = 10'd316;
assign feature_index_9[276] = 10'd354;
assign feature_index_9[277] = 10'd271;
assign feature_index_9[278] = 10'd383;
assign feature_index_9[279] = 10'd215;
assign feature_index_9[280] = 10'd635;
assign feature_index_9[281] = 10'd0;
assign feature_index_9[282] = 10'd0;
assign feature_index_9[283] = 10'd0;
assign feature_index_9[284] = 10'd0;
assign feature_index_9[285] = 10'd0;
assign feature_index_9[286] = 10'd0;
assign feature_index_9[287] = 10'd185;
assign feature_index_9[288] = 10'd622;
assign feature_index_9[289] = 10'd401;
assign feature_index_9[290] = 10'd237;
assign feature_index_9[291] = 10'd514;
assign feature_index_9[292] = 10'd486;
assign feature_index_9[293] = 10'd567;
assign feature_index_9[294] = 10'd135;
assign feature_index_9[295] = 10'd515;
assign feature_index_9[296] = 10'd160;
assign feature_index_9[297] = 10'd623;
assign feature_index_9[298] = 10'd327;
assign feature_index_9[299] = 10'd154;
assign feature_index_9[300] = 10'd457;
assign feature_index_9[301] = 10'd490;
assign feature_index_9[302] = 10'd443;
assign feature_index_9[303] = 10'd468;
assign feature_index_9[304] = 10'd519;
assign feature_index_9[305] = 10'd266;
assign feature_index_9[306] = 10'd100;
assign feature_index_9[307] = 10'd0;
assign feature_index_9[308] = 10'd578;
assign feature_index_9[309] = 10'd0;
assign feature_index_9[310] = 10'd0;
assign feature_index_9[311] = 10'd433;
assign feature_index_9[312] = 10'd627;
assign feature_index_9[313] = 10'd379;
assign feature_index_9[314] = 10'd191;
assign feature_index_9[315] = 10'd519;
assign feature_index_9[316] = 10'd652;
assign feature_index_9[317] = 10'd519;
assign feature_index_9[318] = 10'd352;
assign feature_index_9[319] = 10'd412;
assign feature_index_9[320] = 10'd710;
assign feature_index_9[321] = 10'd379;
assign feature_index_9[322] = 10'd374;
assign feature_index_9[323] = 10'd262;
assign feature_index_9[324] = 10'd0;
assign feature_index_9[325] = 10'd382;
assign feature_index_9[326] = 10'd542;
assign feature_index_9[327] = 10'd514;
assign feature_index_9[328] = 10'd248;
assign feature_index_9[329] = 10'd180;
assign feature_index_9[330] = 10'd602;
assign feature_index_9[331] = 10'd659;
assign feature_index_9[332] = 10'd358;
assign feature_index_9[333] = 10'd569;
assign feature_index_9[334] = 10'd330;
assign feature_index_9[335] = 10'd374;
assign feature_index_9[336] = 10'd408;
assign feature_index_9[337] = 10'd345;
assign feature_index_9[338] = 10'd0;
assign feature_index_9[339] = 10'd543;
assign feature_index_9[340] = 10'd631;
assign feature_index_9[341] = 10'd0;
assign feature_index_9[342] = 10'd317;
assign feature_index_9[343] = 10'd623;
assign feature_index_9[344] = 10'd326;
assign feature_index_9[345] = 10'd594;
assign feature_index_9[346] = 10'd344;
assign feature_index_9[347] = 10'd682;
assign feature_index_9[348] = 10'd0;
assign feature_index_9[349] = 10'd406;
assign feature_index_9[350] = 10'd131;
assign feature_index_9[351] = 10'd407;
assign feature_index_9[352] = 10'd358;
assign feature_index_9[353] = 10'd498;
assign feature_index_9[354] = 10'd480;
assign feature_index_9[355] = 10'd184;
assign feature_index_9[356] = 10'd341;
assign feature_index_9[357] = 10'd0;
assign feature_index_9[358] = 10'd0;
assign feature_index_9[359] = 10'd0;
assign feature_index_9[360] = 10'd240;
assign feature_index_9[361] = 10'd440;
assign feature_index_9[362] = 10'd433;
assign feature_index_9[363] = 10'd664;
assign feature_index_9[364] = 10'd386;
assign feature_index_9[365] = 10'd0;
assign feature_index_9[366] = 10'd578;
assign feature_index_9[367] = 10'd105;
assign feature_index_9[368] = 10'd720;
assign feature_index_9[369] = 10'd577;
assign feature_index_9[370] = 10'd349;
assign feature_index_9[371] = 10'd606;
assign feature_index_9[372] = 10'd154;
assign feature_index_9[373] = 10'd161;
assign feature_index_9[374] = 10'd624;
assign feature_index_9[375] = 10'd488;
assign feature_index_9[376] = 10'd320;
assign feature_index_9[377] = 10'd0;
assign feature_index_9[378] = 10'd0;
assign feature_index_9[379] = 10'd0;
assign feature_index_9[380] = 10'd319;
assign feature_index_9[381] = 10'd536;
assign feature_index_9[382] = 10'd435;
assign feature_index_9[383] = 10'd465;
assign feature_index_9[384] = 10'd403;
assign feature_index_9[385] = 10'd583;
assign feature_index_9[386] = 10'd263;
assign feature_index_9[387] = 10'd317;
assign feature_index_9[388] = 10'd595;
assign feature_index_9[389] = 10'd624;
assign feature_index_9[390] = 10'd185;
assign feature_index_9[391] = 10'd433;
assign feature_index_9[392] = 10'd542;
assign feature_index_9[393] = 10'd374;
assign feature_index_9[394] = 10'd351;
assign feature_index_9[395] = 10'd549;
assign feature_index_9[396] = 10'd545;
assign feature_index_9[397] = 10'd624;
assign feature_index_9[398] = 10'd353;
assign feature_index_9[399] = 10'd740;
assign feature_index_9[400] = 10'd574;
assign feature_index_9[401] = 10'd431;
assign feature_index_9[402] = 10'd0;
assign feature_index_9[403] = 10'd180;
assign feature_index_9[404] = 10'd179;
assign feature_index_9[405] = 10'd602;
assign feature_index_9[406] = 10'd573;
assign feature_index_9[407] = 10'd486;
assign feature_index_9[408] = 10'd543;
assign feature_index_9[409] = 10'd711;
assign feature_index_9[410] = 10'd325;
assign feature_index_9[411] = 10'd159;
assign feature_index_9[412] = 10'd265;
assign feature_index_9[413] = 10'd209;
assign feature_index_9[414] = 10'd543;
assign feature_index_9[415] = 10'd153;
assign feature_index_9[416] = 10'd439;
assign feature_index_9[417] = 10'd0;
assign feature_index_9[418] = 10'd0;
assign feature_index_9[419] = 10'd299;
assign feature_index_9[420] = 10'd0;
assign feature_index_9[421] = 10'd0;
assign feature_index_9[422] = 10'd0;
assign feature_index_9[423] = 10'd377;
assign feature_index_9[424] = 10'd544;
assign feature_index_9[425] = 10'd427;
assign feature_index_9[426] = 10'd517;
assign feature_index_9[427] = 10'd739;
assign feature_index_9[428] = 10'd595;
assign feature_index_9[429] = 10'd0;
assign feature_index_9[430] = 10'd259;
assign feature_index_9[431] = 10'd374;
assign feature_index_9[432] = 10'd0;
assign feature_index_9[433] = 10'd567;
assign feature_index_9[434] = 10'd443;
assign feature_index_9[435] = 10'd315;
assign feature_index_9[436] = 10'd158;
assign feature_index_9[437] = 10'd288;
assign feature_index_9[438] = 10'd548;
assign feature_index_9[439] = 10'd427;
assign feature_index_9[440] = 10'd183;
assign feature_index_9[441] = 10'd570;
assign feature_index_9[442] = 10'd321;
assign feature_index_9[443] = 10'd155;
assign feature_index_9[444] = 10'd0;
assign feature_index_9[445] = 10'd654;
assign feature_index_9[446] = 10'd443;
assign feature_index_9[447] = 10'd403;
assign feature_index_9[448] = 10'd320;
assign feature_index_9[449] = 10'd603;
assign feature_index_9[450] = 10'd0;
assign feature_index_9[451] = 10'd427;
assign feature_index_9[452] = 10'd378;
assign feature_index_9[453] = 10'd483;
assign feature_index_9[454] = 10'd600;
assign feature_index_9[455] = 10'd514;
assign feature_index_9[456] = 10'd319;
assign feature_index_9[457] = 10'd459;
assign feature_index_9[458] = 10'd0;
assign feature_index_9[459] = 10'd92;
assign feature_index_9[460] = 10'd341;
assign feature_index_9[461] = 10'd407;
assign feature_index_9[462] = 10'd540;
assign feature_index_9[463] = 10'd654;
assign feature_index_9[464] = 10'd690;
assign feature_index_9[465] = 10'd708;
assign feature_index_9[466] = 10'd663;
assign feature_index_9[467] = 10'd179;
assign feature_index_9[468] = 10'd372;
assign feature_index_9[469] = 10'd544;
assign feature_index_9[470] = 10'd485;
assign feature_index_9[471] = 10'd217;
assign feature_index_9[472] = 10'd543;
assign feature_index_9[473] = 10'd651;
assign feature_index_9[474] = 10'd487;
assign feature_index_9[475] = 10'd375;
assign feature_index_9[476] = 10'd0;
assign feature_index_9[477] = 10'd399;
assign feature_index_9[478] = 10'd428;
assign feature_index_9[479] = 10'd323;
assign feature_index_9[480] = 10'd0;
assign feature_index_9[481] = 10'd239;
assign feature_index_9[482] = 10'd236;
assign feature_index_9[483] = 10'd469;
assign feature_index_9[484] = 10'd272;
assign feature_index_9[485] = 10'd355;
assign feature_index_9[486] = 10'd159;
assign feature_index_9[487] = 10'd243;
assign feature_index_9[488] = 10'd290;
assign feature_index_9[489] = 10'd261;
assign feature_index_9[490] = 10'd567;
assign feature_index_9[491] = 10'd379;
assign feature_index_9[492] = 10'd292;
assign feature_index_9[493] = 10'd658;
assign feature_index_9[494] = 10'd658;
assign feature_index_9[495] = 10'd376;
assign feature_index_9[496] = 10'd297;
assign feature_index_9[497] = 10'd401;
assign feature_index_9[498] = 10'd403;
assign feature_index_9[499] = 10'd511;
assign feature_index_9[500] = 10'd412;
assign feature_index_9[501] = 10'd538;
assign feature_index_9[502] = 10'd453;
assign feature_index_9[503] = 10'd349;
assign feature_index_9[504] = 10'd102;
assign feature_index_9[505] = 10'd628;
assign feature_index_9[506] = 10'd295;
assign feature_index_9[507] = 10'd0;
assign feature_index_9[508] = 10'd544;
assign feature_index_9[509] = 10'd377;
assign feature_index_9[510] = 10'd426;
assign feature_index_9[511] = 10'd685;
assign feature_index_9[512] = 10'd132;
assign feature_index_9[513] = 10'd303;
assign feature_index_9[514] = 10'd384;
assign feature_index_9[515] = 10'd374;
assign feature_index_9[516] = 10'd105;
assign feature_index_9[517] = 10'd545;
assign feature_index_9[518] = 10'd622;
assign feature_index_9[519] = 10'd383;
assign feature_index_9[520] = 10'd184;
assign feature_index_9[521] = 10'd0;
assign feature_index_9[522] = 10'd0;
assign feature_index_9[523] = 10'd213;
assign feature_index_9[524] = 10'd182;
assign feature_index_9[525] = 10'd0;
assign feature_index_9[526] = 10'd429;
assign feature_index_9[527] = 10'd211;
assign feature_index_9[528] = 10'd577;
assign feature_index_9[529] = 10'd351;
assign feature_index_9[530] = 10'd378;
assign feature_index_9[531] = 10'd572;
assign feature_index_9[532] = 10'd572;
assign feature_index_9[533] = 10'd372;
assign feature_index_9[534] = 10'd270;
assign feature_index_9[535] = 10'd178;
assign feature_index_9[536] = 10'd543;
assign feature_index_9[537] = 10'd211;
assign feature_index_9[538] = 10'd154;
assign feature_index_9[539] = 10'd377;
assign feature_index_9[540] = 10'd262;
assign feature_index_9[541] = 10'd341;
assign feature_index_9[542] = 10'd556;
assign feature_index_9[543] = 10'd298;
assign feature_index_9[544] = 10'd0;
assign feature_index_9[545] = 10'd0;
assign feature_index_9[546] = 10'd0;
assign feature_index_9[547] = 10'd0;
assign feature_index_9[548] = 10'd0;
assign feature_index_9[549] = 10'd0;
assign feature_index_9[550] = 10'd0;
assign feature_index_9[551] = 10'd0;
assign feature_index_9[552] = 10'd347;
assign feature_index_9[553] = 10'd322;
assign feature_index_9[554] = 10'd689;
assign feature_index_9[555] = 10'd0;
assign feature_index_9[556] = 10'd0;
assign feature_index_9[557] = 10'd0;
assign feature_index_9[558] = 10'd242;
assign feature_index_9[559] = 10'd229;
assign feature_index_9[560] = 10'd0;
assign feature_index_9[561] = 10'd351;
assign feature_index_9[562] = 10'd324;
assign feature_index_9[563] = 10'd0;
assign feature_index_9[564] = 10'd0;
assign feature_index_9[565] = 10'd0;
assign feature_index_9[566] = 10'd0;
assign feature_index_9[567] = 10'd0;
assign feature_index_9[568] = 10'd0;
assign feature_index_9[569] = 10'd0;
assign feature_index_9[570] = 10'd0;
assign feature_index_9[571] = 10'd0;
assign feature_index_9[572] = 10'd0;
assign feature_index_9[573] = 10'd0;
assign feature_index_9[574] = 10'd0;
assign feature_index_9[575] = 10'd685;
assign feature_index_9[576] = 10'd122;
assign feature_index_9[577] = 10'd161;
assign feature_index_9[578] = 10'd355;
assign feature_index_9[579] = 10'd234;
assign feature_index_9[580] = 10'd549;
assign feature_index_9[581] = 10'd592;
assign feature_index_9[582] = 10'd374;
assign feature_index_9[583] = 10'd263;
assign feature_index_9[584] = 10'd439;
assign feature_index_9[585] = 10'd291;
assign feature_index_9[586] = 10'd321;
assign feature_index_9[587] = 10'd352;
assign feature_index_9[588] = 10'd0;
assign feature_index_9[589] = 10'd497;
assign feature_index_9[590] = 10'd522;
assign feature_index_9[591] = 10'd163;
assign feature_index_9[592] = 10'd270;
assign feature_index_9[593] = 10'd426;
assign feature_index_9[594] = 10'd265;
assign feature_index_9[595] = 10'd265;
assign feature_index_9[596] = 10'd162;
assign feature_index_9[597] = 10'd653;
assign feature_index_9[598] = 10'd598;
assign feature_index_9[599] = 10'd464;
assign feature_index_9[600] = 10'd212;
assign feature_index_9[601] = 10'd411;
assign feature_index_9[602] = 10'd495;
assign feature_index_9[603] = 10'd609;
assign feature_index_9[604] = 10'd319;
assign feature_index_9[605] = 10'd0;
assign feature_index_9[606] = 10'd567;
assign feature_index_9[607] = 10'd460;
assign feature_index_9[608] = 10'd241;
assign feature_index_9[609] = 10'd325;
assign feature_index_9[610] = 10'd429;
assign feature_index_9[611] = 10'd513;
assign feature_index_9[612] = 10'd150;
assign feature_index_9[613] = 10'd296;
assign feature_index_9[614] = 10'd243;
assign feature_index_9[615] = 10'd0;
assign feature_index_9[616] = 10'd0;
assign feature_index_9[617] = 10'd0;
assign feature_index_9[618] = 10'd0;
assign feature_index_9[619] = 10'd0;
assign feature_index_9[620] = 10'd0;
assign feature_index_9[621] = 10'd0;
assign feature_index_9[622] = 10'd0;
assign feature_index_9[623] = 10'd0;
assign feature_index_9[624] = 10'd0;
assign feature_index_9[625] = 10'd259;
assign feature_index_9[626] = 10'd0;
assign feature_index_9[627] = 10'd376;
assign feature_index_9[628] = 10'd385;
assign feature_index_9[629] = 10'd216;
assign feature_index_9[630] = 10'd0;
assign feature_index_9[631] = 10'd0;
assign feature_index_9[632] = 10'd215;
assign feature_index_9[633] = 10'd287;
assign feature_index_9[634] = 10'd496;
assign feature_index_9[635] = 10'd0;
assign feature_index_9[636] = 10'd0;
assign feature_index_9[637] = 10'd549;
assign feature_index_9[638] = 10'd294;
assign feature_index_9[639] = 10'd354;
assign feature_index_9[640] = 10'd372;
assign feature_index_9[641] = 10'd416;
assign feature_index_9[642] = 10'd0;
assign feature_index_9[643] = 10'd494;
assign feature_index_9[644] = 10'd217;
assign feature_index_9[645] = 10'd512;
assign feature_index_9[646] = 10'd739;
assign feature_index_9[647] = 10'd370;
assign feature_index_9[648] = 10'd0;
assign feature_index_9[649] = 10'd0;
assign feature_index_9[650] = 10'd0;
assign feature_index_9[651] = 10'd461;
assign feature_index_9[652] = 10'd508;
assign feature_index_9[653] = 10'd0;
assign feature_index_9[654] = 10'd0;
assign feature_index_9[655] = 10'd270;
assign feature_index_9[656] = 10'd595;
assign feature_index_9[657] = 10'd237;
assign feature_index_9[658] = 10'd357;
assign feature_index_9[659] = 10'd0;
assign feature_index_9[660] = 10'd491;
assign feature_index_9[661] = 10'd0;
assign feature_index_9[662] = 10'd608;
assign feature_index_9[663] = 10'd240;
assign feature_index_9[664] = 10'd212;
assign feature_index_9[665] = 10'd0;
assign feature_index_9[666] = 10'd0;
assign feature_index_9[667] = 10'd241;
assign feature_index_9[668] = 10'd212;
assign feature_index_9[669] = 10'd566;
assign feature_index_9[670] = 10'd383;
assign feature_index_9[671] = 10'd683;
assign feature_index_9[672] = 10'd175;
assign feature_index_9[673] = 10'd497;
assign feature_index_9[674] = 10'd344;
assign feature_index_9[675] = 10'd0;
assign feature_index_9[676] = 10'd0;
assign feature_index_9[677] = 10'd0;
assign feature_index_9[678] = 10'd0;
assign feature_index_9[679] = 10'd175;
assign feature_index_9[680] = 10'd246;
assign feature_index_9[681] = 10'd0;
assign feature_index_9[682] = 10'd327;
assign feature_index_9[683] = 10'd0;
assign feature_index_9[684] = 10'd0;
assign feature_index_9[685] = 10'd0;
assign feature_index_9[686] = 10'd630;
assign feature_index_9[687] = 10'd459;
assign feature_index_9[688] = 10'd593;
assign feature_index_9[689] = 10'd598;
assign feature_index_9[690] = 10'd680;
assign feature_index_9[691] = 10'd345;
assign feature_index_9[692] = 10'd630;
assign feature_index_9[693] = 10'd330;
assign feature_index_9[694] = 10'd440;
assign feature_index_9[695] = 10'd160;
assign feature_index_9[696] = 10'd567;
assign feature_index_9[697] = 10'd0;
assign feature_index_9[698] = 10'd0;
assign feature_index_9[699] = 10'd288;
assign feature_index_9[700] = 10'd592;
assign feature_index_9[701] = 10'd230;
assign feature_index_9[702] = 10'd0;
assign feature_index_9[703] = 10'd598;
assign feature_index_9[704] = 10'd331;
assign feature_index_9[705] = 10'd384;
assign feature_index_9[706] = 10'd236;
assign feature_index_9[707] = 10'd266;
assign feature_index_9[708] = 10'd410;
assign feature_index_9[709] = 10'd438;
assign feature_index_9[710] = 10'd547;
assign feature_index_9[711] = 10'd495;
assign feature_index_9[712] = 10'd162;
assign feature_index_9[713] = 10'd683;
assign feature_index_9[714] = 10'd0;
assign feature_index_9[715] = 10'd0;
assign feature_index_9[716] = 10'd0;
assign feature_index_9[717] = 10'd0;
assign feature_index_9[718] = 10'd0;
assign feature_index_9[719] = 10'd0;
assign feature_index_9[720] = 10'd0;
assign feature_index_9[721] = 10'd130;
assign feature_index_9[722] = 10'd553;
assign feature_index_9[723] = 10'd0;
assign feature_index_9[724] = 10'd0;
assign feature_index_9[725] = 10'd465;
assign feature_index_9[726] = 10'd0;
assign feature_index_9[727] = 10'd0;
assign feature_index_9[728] = 10'd322;
assign feature_index_9[729] = 10'd440;
assign feature_index_9[730] = 10'd429;
assign feature_index_9[731] = 10'd0;
assign feature_index_9[732] = 10'd0;
assign feature_index_9[733] = 10'd0;
assign feature_index_9[734] = 10'd0;
assign feature_index_9[735] = 10'd597;
assign feature_index_9[736] = 10'd0;
assign feature_index_9[737] = 10'd241;
assign feature_index_9[738] = 10'd289;
assign feature_index_9[739] = 10'd434;
assign feature_index_9[740] = 10'd239;
assign feature_index_9[741] = 10'd0;
assign feature_index_9[742] = 10'd351;
assign feature_index_9[743] = 10'd597;
assign feature_index_9[744] = 10'd604;
assign feature_index_9[745] = 10'd0;
assign feature_index_9[746] = 10'd331;
assign feature_index_9[747] = 10'd0;
assign feature_index_9[748] = 10'd0;
assign feature_index_9[749] = 10'd570;
assign feature_index_9[750] = 10'd343;
assign feature_index_9[751] = 10'd432;
assign feature_index_9[752] = 10'd346;
assign feature_index_9[753] = 10'd211;
assign feature_index_9[754] = 10'd176;
assign feature_index_9[755] = 10'd0;
assign feature_index_9[756] = 10'd0;
assign feature_index_9[757] = 10'd0;
assign feature_index_9[758] = 10'd0;
assign feature_index_9[759] = 10'd0;
assign feature_index_9[760] = 10'd0;
assign feature_index_9[761] = 10'd490;
assign feature_index_9[762] = 10'd522;
assign feature_index_9[763] = 10'd547;
assign feature_index_9[764] = 10'd128;
assign feature_index_9[765] = 10'd410;
assign feature_index_9[766] = 10'd540;
assign feature_index_9[767] = 10'd430;
assign feature_index_9[768] = 10'd490;
assign feature_index_9[769] = 10'd157;
assign feature_index_9[770] = 10'd157;
assign feature_index_9[771] = 10'd466;
assign feature_index_9[772] = 10'd187;
assign feature_index_9[773] = 10'd433;
assign feature_index_9[774] = 10'd524;
assign feature_index_9[775] = 10'd657;
assign feature_index_9[776] = 10'd175;
assign feature_index_9[777] = 10'd235;
assign feature_index_9[778] = 10'd493;
assign feature_index_9[779] = 10'd150;
assign feature_index_9[780] = 10'd292;
assign feature_index_9[781] = 10'd267;
assign feature_index_9[782] = 10'd377;
assign feature_index_9[783] = 10'd156;
assign feature_index_9[784] = 10'd230;
assign feature_index_9[785] = 10'd154;
assign feature_index_9[786] = 10'd605;
assign feature_index_9[787] = 10'd399;
assign feature_index_9[788] = 10'd323;
assign feature_index_9[789] = 10'd266;
assign feature_index_9[790] = 10'd0;
assign feature_index_9[791] = 10'd652;
assign feature_index_9[792] = 10'd325;
assign feature_index_9[793] = 10'd316;
assign feature_index_9[794] = 10'd262;
assign feature_index_9[795] = 10'd320;
assign feature_index_9[796] = 10'd460;
assign feature_index_9[797] = 10'd0;
assign feature_index_9[798] = 10'd0;
assign feature_index_9[799] = 10'd210;
assign feature_index_9[800] = 10'd402;
assign feature_index_9[801] = 10'd327;
assign feature_index_9[802] = 10'd343;
assign feature_index_9[803] = 10'd350;
assign feature_index_9[804] = 10'd95;
assign feature_index_9[805] = 10'd0;
assign feature_index_9[806] = 10'd0;
assign feature_index_9[807] = 10'd458;
assign feature_index_9[808] = 10'd321;
assign feature_index_9[809] = 10'd552;
assign feature_index_9[810] = 10'd343;
assign feature_index_9[811] = 10'd633;
assign feature_index_9[812] = 10'd379;
assign feature_index_9[813] = 10'd292;
assign feature_index_9[814] = 10'd317;
assign feature_index_9[815] = 10'd188;
assign feature_index_9[816] = 10'd322;
assign feature_index_9[817] = 10'd594;
assign feature_index_9[818] = 10'd99;
assign feature_index_9[819] = 10'd624;
assign feature_index_9[820] = 10'd295;
assign feature_index_9[821] = 10'd659;
assign feature_index_9[822] = 10'd658;
assign feature_index_9[823] = 10'd203;
assign feature_index_9[824] = 10'd602;
assign feature_index_9[825] = 10'd656;
assign feature_index_9[826] = 10'd215;
assign feature_index_9[827] = 10'd296;
assign feature_index_9[828] = 10'd716;
assign feature_index_9[829] = 10'd190;
assign feature_index_9[830] = 10'd412;
assign feature_index_9[831] = 10'd93;
assign feature_index_9[832] = 10'd155;
assign feature_index_9[833] = 10'd464;
assign feature_index_9[834] = 10'd235;
assign feature_index_9[835] = 10'd0;
assign feature_index_9[836] = 10'd0;
assign feature_index_9[837] = 10'd0;
assign feature_index_9[838] = 10'd0;
assign feature_index_9[839] = 10'd0;
assign feature_index_9[840] = 10'd516;
assign feature_index_9[841] = 10'd0;
assign feature_index_9[842] = 10'd0;
assign feature_index_9[843] = 10'd0;
assign feature_index_9[844] = 10'd0;
assign feature_index_9[845] = 10'd0;
assign feature_index_9[846] = 10'd0;
assign feature_index_9[847] = 10'd0;
assign feature_index_9[848] = 10'd0;
assign feature_index_9[849] = 10'd353;
assign feature_index_9[850] = 10'd0;
assign feature_index_9[851] = 10'd0;
assign feature_index_9[852] = 10'd469;
assign feature_index_9[853] = 10'd368;
assign feature_index_9[854] = 10'd598;
assign feature_index_9[855] = 10'd322;
assign feature_index_9[856] = 10'd330;
assign feature_index_9[857] = 10'd468;
assign feature_index_9[858] = 10'd0;
assign feature_index_9[859] = 10'd0;
assign feature_index_9[860] = 10'd0;
assign feature_index_9[861] = 10'd0;
assign feature_index_9[862] = 10'd0;
assign feature_index_9[863] = 10'd354;
assign feature_index_9[864] = 10'd474;
assign feature_index_9[865] = 10'd0;
assign feature_index_9[866] = 10'd0;
assign feature_index_9[867] = 10'd443;
assign feature_index_9[868] = 10'd177;
assign feature_index_9[869] = 10'd289;
assign feature_index_9[870] = 10'd686;
assign feature_index_9[871] = 10'd455;
assign feature_index_9[872] = 10'd516;
assign feature_index_9[873] = 10'd125;
assign feature_index_9[874] = 10'd177;
assign feature_index_9[875] = 10'd483;
assign feature_index_9[876] = 10'd469;
assign feature_index_9[877] = 10'd325;
assign feature_index_9[878] = 10'd191;
assign feature_index_9[879] = 10'd97;
assign feature_index_9[880] = 10'd744;
assign feature_index_9[881] = 10'd128;
assign feature_index_9[882] = 10'd321;
assign feature_index_9[883] = 10'd544;
assign feature_index_9[884] = 10'd212;
assign feature_index_9[885] = 10'd300;
assign feature_index_9[886] = 10'd0;
assign feature_index_9[887] = 10'd189;
assign feature_index_9[888] = 10'd523;
assign feature_index_9[889] = 10'd0;
assign feature_index_9[890] = 10'd0;
assign feature_index_9[891] = 10'd258;
assign feature_index_9[892] = 10'd351;
assign feature_index_9[893] = 10'd0;
assign feature_index_9[894] = 10'd147;
assign feature_index_9[895] = 10'd467;
assign feature_index_9[896] = 10'd130;
assign feature_index_9[897] = 10'd265;
assign feature_index_9[898] = 10'd574;
assign feature_index_9[899] = 10'd625;
assign feature_index_9[900] = 10'd655;
assign feature_index_9[901] = 10'd0;
assign feature_index_9[902] = 10'd0;
assign feature_index_9[903] = 10'd264;
assign feature_index_9[904] = 10'd424;
assign feature_index_9[905] = 10'd603;
assign feature_index_9[906] = 10'd510;
assign feature_index_9[907] = 10'd300;
assign feature_index_9[908] = 10'd288;
assign feature_index_9[909] = 10'd345;
assign feature_index_9[910] = 10'd271;
assign feature_index_9[911] = 10'd0;
assign feature_index_9[912] = 10'd162;
assign feature_index_9[913] = 10'd241;
assign feature_index_9[914] = 10'd0;
assign feature_index_9[915] = 10'd405;
assign feature_index_9[916] = 10'd348;
assign feature_index_9[917] = 10'd0;
assign feature_index_9[918] = 10'd0;
assign feature_index_9[919] = 10'd295;
assign feature_index_9[920] = 10'd0;
assign feature_index_9[921] = 10'd627;
assign feature_index_9[922] = 10'd0;
assign feature_index_9[923] = 10'd0;
assign feature_index_9[924] = 10'd706;
assign feature_index_9[925] = 10'd400;
assign feature_index_9[926] = 10'd325;
assign feature_index_9[927] = 10'd179;
assign feature_index_9[928] = 10'd682;
assign feature_index_9[929] = 10'd566;
assign feature_index_9[930] = 10'd0;
assign feature_index_9[931] = 10'd181;
assign feature_index_9[932] = 10'd359;
assign feature_index_9[933] = 10'd626;
assign feature_index_9[934] = 10'd230;
assign feature_index_9[935] = 10'd635;
assign feature_index_9[936] = 10'd316;
assign feature_index_9[937] = 10'd542;
assign feature_index_9[938] = 10'd353;
assign feature_index_9[939] = 10'd515;
assign feature_index_9[940] = 10'd332;
assign feature_index_9[941] = 10'd287;
assign feature_index_9[942] = 10'd343;
assign feature_index_9[943] = 10'd242;
assign feature_index_9[944] = 10'd486;
assign feature_index_9[945] = 10'd515;
assign feature_index_9[946] = 10'd488;
assign feature_index_9[947] = 10'd276;
assign feature_index_9[948] = 10'd496;
assign feature_index_9[949] = 10'd329;
assign feature_index_9[950] = 10'd130;
assign feature_index_9[951] = 10'd665;
assign feature_index_9[952] = 10'd292;
assign feature_index_9[953] = 10'd0;
assign feature_index_9[954] = 10'd0;
assign feature_index_9[955] = 10'd486;
assign feature_index_9[956] = 10'd602;
assign feature_index_9[957] = 10'd459;
assign feature_index_9[958] = 10'd304;
assign feature_index_9[959] = 10'd546;
assign feature_index_9[960] = 10'd460;
assign feature_index_9[961] = 10'd0;
assign feature_index_9[962] = 10'd0;
assign feature_index_9[963] = 10'd238;
assign feature_index_9[964] = 10'd436;
assign feature_index_9[965] = 10'd0;
assign feature_index_9[966] = 10'd628;
assign feature_index_9[967] = 10'd289;
assign feature_index_9[968] = 10'd247;
assign feature_index_9[969] = 10'd347;
assign feature_index_9[970] = 10'd518;
assign feature_index_9[971] = 10'd465;
assign feature_index_9[972] = 10'd206;
assign feature_index_9[973] = 10'd0;
assign feature_index_9[974] = 10'd0;
assign feature_index_9[975] = 10'd296;
assign feature_index_9[976] = 10'd326;
assign feature_index_9[977] = 10'd375;
assign feature_index_9[978] = 10'd496;
assign feature_index_9[979] = 10'd606;
assign feature_index_9[980] = 10'd405;
assign feature_index_9[981] = 10'd244;
assign feature_index_9[982] = 10'd316;
assign feature_index_9[983] = 10'd333;
assign feature_index_9[984] = 10'd377;
assign feature_index_9[985] = 10'd301;
assign feature_index_9[986] = 10'd630;
assign feature_index_9[987] = 10'd380;
assign feature_index_9[988] = 10'd520;
assign feature_index_9[989] = 10'd191;
assign feature_index_9[990] = 10'd387;
assign feature_index_9[991] = 10'd434;
assign feature_index_9[992] = 10'd601;
assign feature_index_9[993] = 10'd0;
assign feature_index_9[994] = 10'd174;
assign feature_index_9[995] = 10'd467;
assign feature_index_9[996] = 10'd158;
assign feature_index_9[997] = 10'd376;
assign feature_index_9[998] = 10'd593;
assign feature_index_9[999] = 10'd544;
assign feature_index_9[1000] = 10'd547;
assign feature_index_9[1001] = 10'd572;
assign feature_index_9[1002] = 10'd159;
assign feature_index_9[1003] = 10'd626;
assign feature_index_9[1004] = 10'd631;
assign feature_index_9[1005] = 10'd436;
assign feature_index_9[1006] = 10'd605;
assign feature_index_9[1007] = 10'd0;
assign feature_index_9[1008] = 10'd0;
assign feature_index_9[1009] = 10'd0;
assign feature_index_9[1010] = 10'd521;
assign feature_index_9[1011] = 10'd0;
assign feature_index_9[1012] = 10'd405;
assign feature_index_9[1013] = 10'd323;
assign feature_index_9[1014] = 10'd466;
assign feature_index_9[1015] = 10'd0;
assign feature_index_9[1016] = 10'd0;
assign feature_index_9[1017] = 10'd325;
assign feature_index_9[1018] = 10'd325;
assign feature_index_9[1019] = 10'd321;
assign feature_index_9[1020] = 10'd494;
assign feature_index_9[1021] = 10'd406;
assign feature_index_9[1022] = 10'd314;

endmodule
